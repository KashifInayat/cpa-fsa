module Mesh( // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177051.2]
  input         clock, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177052.4]
  input  [7:0]  io_in_a_0_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input  [7:0]  io_in_a_1_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input  [7:0]  io_in_a_2_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input  [7:0]  io_in_a_3_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input  [7:0]  io_in_a_4_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input  [7:0]  io_in_a_5_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input  [7:0]  io_in_a_6_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input  [7:0]  io_in_a_7_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input  [7:0]  io_in_d_0_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input  [7:0]  io_in_d_1_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input  [7:0]  io_in_d_2_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input  [7:0]  io_in_d_3_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input  [7:0]  io_in_d_4_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input  [7:0]  io_in_d_5_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input  [7:0]  io_in_d_6_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input  [7:0]  io_in_d_7_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input  [7:0]  io_in_b_0_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input  [7:0]  io_in_b_1_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input  [7:0]  io_in_b_2_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input  [7:0]  io_in_b_3_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input  [7:0]  io_in_b_4_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input  [7:0]  io_in_b_5_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input  [7:0]  io_in_b_6_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input  [7:0]  io_in_b_7_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input         io_in_control_0_0_propagate, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input  [4:0]  io_in_control_0_0_shift, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input         io_in_control_1_0_propagate, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input  [4:0]  io_in_control_1_0_shift, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input         io_in_control_2_0_propagate, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input  [4:0]  io_in_control_2_0_shift, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input         io_in_control_3_0_propagate, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input  [4:0]  io_in_control_3_0_shift, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input         io_in_control_4_0_propagate, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input  [4:0]  io_in_control_4_0_shift, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input         io_in_control_5_0_propagate, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input  [4:0]  io_in_control_5_0_shift, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input         io_in_control_6_0_propagate, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input  [4:0]  io_in_control_6_0_shift, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input         io_in_control_7_0_propagate, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input  [4:0]  io_in_control_7_0_shift, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  output [18:0] io_out_c_0_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  output [18:0] io_out_c_1_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  output [18:0] io_out_c_2_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  output [18:0] io_out_c_3_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  output [18:0] io_out_c_4_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  output [18:0] io_out_c_5_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  output [18:0] io_out_c_6_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  output [18:0] io_out_c_7_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  output [18:0] io_out_b_0_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  output [18:0] io_out_b_1_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  output [18:0] io_out_b_2_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  output [18:0] io_out_b_3_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  output [18:0] io_out_b_4_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  output [18:0] io_out_b_5_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  output [18:0] io_out_b_6_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  output [18:0] io_out_b_7_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input         io_in_valid_0_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input         io_in_valid_1_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input         io_in_valid_2_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input         io_in_valid_3_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input         io_in_valid_4_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input         io_in_valid_5_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input         io_in_valid_6_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  input         io_in_valid_7_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
  output        io_out_valid_0_0 // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177054.4]
);
  wire  mesh_0_0_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177056.4]
  wire [7:0] mesh_0_0_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177056.4]
  wire [18:0] mesh_0_0_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177056.4]
  wire [18:0] mesh_0_0_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177056.4]
  wire  mesh_0_0_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177056.4]
  wire [4:0] mesh_0_0_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177056.4]
  wire [7:0] mesh_0_0_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177056.4]
  wire [18:0] mesh_0_0_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177056.4]
  wire [18:0] mesh_0_0_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177056.4]
  wire  mesh_0_0_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177056.4]
  wire [4:0] mesh_0_0_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177056.4]
  wire  mesh_0_0_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177056.4]
  wire  mesh_0_0_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177056.4]
  wire  mesh_0_1_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177059.4]
  wire [7:0] mesh_0_1_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177059.4]
  wire [18:0] mesh_0_1_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177059.4]
  wire [18:0] mesh_0_1_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177059.4]
  wire  mesh_0_1_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177059.4]
  wire [4:0] mesh_0_1_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177059.4]
  wire [7:0] mesh_0_1_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177059.4]
  wire [18:0] mesh_0_1_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177059.4]
  wire [18:0] mesh_0_1_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177059.4]
  wire  mesh_0_1_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177059.4]
  wire [4:0] mesh_0_1_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177059.4]
  wire  mesh_0_1_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177059.4]
  wire  mesh_0_1_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177059.4]
  wire  mesh_0_2_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177062.4]
  wire [7:0] mesh_0_2_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177062.4]
  wire [18:0] mesh_0_2_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177062.4]
  wire [18:0] mesh_0_2_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177062.4]
  wire  mesh_0_2_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177062.4]
  wire [4:0] mesh_0_2_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177062.4]
  wire [7:0] mesh_0_2_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177062.4]
  wire [18:0] mesh_0_2_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177062.4]
  wire [18:0] mesh_0_2_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177062.4]
  wire  mesh_0_2_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177062.4]
  wire [4:0] mesh_0_2_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177062.4]
  wire  mesh_0_2_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177062.4]
  wire  mesh_0_2_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177062.4]
  wire  mesh_0_3_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177065.4]
  wire [7:0] mesh_0_3_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177065.4]
  wire [18:0] mesh_0_3_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177065.4]
  wire [18:0] mesh_0_3_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177065.4]
  wire  mesh_0_3_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177065.4]
  wire [4:0] mesh_0_3_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177065.4]
  wire [7:0] mesh_0_3_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177065.4]
  wire [18:0] mesh_0_3_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177065.4]
  wire [18:0] mesh_0_3_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177065.4]
  wire  mesh_0_3_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177065.4]
  wire [4:0] mesh_0_3_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177065.4]
  wire  mesh_0_3_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177065.4]
  wire  mesh_0_3_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177065.4]
  wire  mesh_0_4_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177068.4]
  wire [7:0] mesh_0_4_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177068.4]
  wire [18:0] mesh_0_4_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177068.4]
  wire [18:0] mesh_0_4_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177068.4]
  wire  mesh_0_4_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177068.4]
  wire [4:0] mesh_0_4_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177068.4]
  wire [7:0] mesh_0_4_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177068.4]
  wire [18:0] mesh_0_4_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177068.4]
  wire [18:0] mesh_0_4_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177068.4]
  wire  mesh_0_4_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177068.4]
  wire [4:0] mesh_0_4_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177068.4]
  wire  mesh_0_4_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177068.4]
  wire  mesh_0_4_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177068.4]
  wire  mesh_0_5_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177071.4]
  wire [7:0] mesh_0_5_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177071.4]
  wire [18:0] mesh_0_5_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177071.4]
  wire [18:0] mesh_0_5_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177071.4]
  wire  mesh_0_5_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177071.4]
  wire [4:0] mesh_0_5_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177071.4]
  wire [7:0] mesh_0_5_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177071.4]
  wire [18:0] mesh_0_5_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177071.4]
  wire [18:0] mesh_0_5_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177071.4]
  wire  mesh_0_5_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177071.4]
  wire [4:0] mesh_0_5_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177071.4]
  wire  mesh_0_5_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177071.4]
  wire  mesh_0_5_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177071.4]
  wire  mesh_0_6_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177074.4]
  wire [7:0] mesh_0_6_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177074.4]
  wire [18:0] mesh_0_6_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177074.4]
  wire [18:0] mesh_0_6_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177074.4]
  wire  mesh_0_6_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177074.4]
  wire [4:0] mesh_0_6_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177074.4]
  wire [7:0] mesh_0_6_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177074.4]
  wire [18:0] mesh_0_6_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177074.4]
  wire [18:0] mesh_0_6_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177074.4]
  wire  mesh_0_6_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177074.4]
  wire [4:0] mesh_0_6_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177074.4]
  wire  mesh_0_6_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177074.4]
  wire  mesh_0_6_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177074.4]
  wire  mesh_0_7_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177077.4]
  wire [7:0] mesh_0_7_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177077.4]
  wire [18:0] mesh_0_7_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177077.4]
  wire [18:0] mesh_0_7_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177077.4]
  wire  mesh_0_7_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177077.4]
  wire [4:0] mesh_0_7_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177077.4]
  wire [7:0] mesh_0_7_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177077.4]
  wire [18:0] mesh_0_7_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177077.4]
  wire [18:0] mesh_0_7_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177077.4]
  wire  mesh_0_7_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177077.4]
  wire [4:0] mesh_0_7_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177077.4]
  wire  mesh_0_7_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177077.4]
  wire  mesh_0_7_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177077.4]
  wire  mesh_1_0_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177080.4]
  wire [7:0] mesh_1_0_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177080.4]
  wire [18:0] mesh_1_0_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177080.4]
  wire [18:0] mesh_1_0_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177080.4]
  wire  mesh_1_0_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177080.4]
  wire [4:0] mesh_1_0_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177080.4]
  wire [7:0] mesh_1_0_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177080.4]
  wire [18:0] mesh_1_0_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177080.4]
  wire [18:0] mesh_1_0_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177080.4]
  wire  mesh_1_0_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177080.4]
  wire [4:0] mesh_1_0_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177080.4]
  wire  mesh_1_0_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177080.4]
  wire  mesh_1_0_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177080.4]
  wire  mesh_1_1_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177083.4]
  wire [7:0] mesh_1_1_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177083.4]
  wire [18:0] mesh_1_1_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177083.4]
  wire [18:0] mesh_1_1_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177083.4]
  wire  mesh_1_1_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177083.4]
  wire [4:0] mesh_1_1_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177083.4]
  wire [7:0] mesh_1_1_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177083.4]
  wire [18:0] mesh_1_1_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177083.4]
  wire [18:0] mesh_1_1_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177083.4]
  wire  mesh_1_1_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177083.4]
  wire [4:0] mesh_1_1_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177083.4]
  wire  mesh_1_1_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177083.4]
  wire  mesh_1_1_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177083.4]
  wire  mesh_1_2_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177086.4]
  wire [7:0] mesh_1_2_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177086.4]
  wire [18:0] mesh_1_2_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177086.4]
  wire [18:0] mesh_1_2_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177086.4]
  wire  mesh_1_2_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177086.4]
  wire [4:0] mesh_1_2_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177086.4]
  wire [7:0] mesh_1_2_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177086.4]
  wire [18:0] mesh_1_2_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177086.4]
  wire [18:0] mesh_1_2_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177086.4]
  wire  mesh_1_2_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177086.4]
  wire [4:0] mesh_1_2_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177086.4]
  wire  mesh_1_2_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177086.4]
  wire  mesh_1_2_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177086.4]
  wire  mesh_1_3_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177089.4]
  wire [7:0] mesh_1_3_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177089.4]
  wire [18:0] mesh_1_3_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177089.4]
  wire [18:0] mesh_1_3_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177089.4]
  wire  mesh_1_3_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177089.4]
  wire [4:0] mesh_1_3_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177089.4]
  wire [7:0] mesh_1_3_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177089.4]
  wire [18:0] mesh_1_3_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177089.4]
  wire [18:0] mesh_1_3_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177089.4]
  wire  mesh_1_3_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177089.4]
  wire [4:0] mesh_1_3_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177089.4]
  wire  mesh_1_3_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177089.4]
  wire  mesh_1_3_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177089.4]
  wire  mesh_1_4_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177092.4]
  wire [7:0] mesh_1_4_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177092.4]
  wire [18:0] mesh_1_4_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177092.4]
  wire [18:0] mesh_1_4_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177092.4]
  wire  mesh_1_4_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177092.4]
  wire [4:0] mesh_1_4_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177092.4]
  wire [7:0] mesh_1_4_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177092.4]
  wire [18:0] mesh_1_4_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177092.4]
  wire [18:0] mesh_1_4_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177092.4]
  wire  mesh_1_4_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177092.4]
  wire [4:0] mesh_1_4_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177092.4]
  wire  mesh_1_4_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177092.4]
  wire  mesh_1_4_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177092.4]
  wire  mesh_1_5_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177095.4]
  wire [7:0] mesh_1_5_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177095.4]
  wire [18:0] mesh_1_5_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177095.4]
  wire [18:0] mesh_1_5_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177095.4]
  wire  mesh_1_5_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177095.4]
  wire [4:0] mesh_1_5_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177095.4]
  wire [7:0] mesh_1_5_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177095.4]
  wire [18:0] mesh_1_5_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177095.4]
  wire [18:0] mesh_1_5_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177095.4]
  wire  mesh_1_5_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177095.4]
  wire [4:0] mesh_1_5_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177095.4]
  wire  mesh_1_5_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177095.4]
  wire  mesh_1_5_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177095.4]
  wire  mesh_1_6_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177098.4]
  wire [7:0] mesh_1_6_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177098.4]
  wire [18:0] mesh_1_6_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177098.4]
  wire [18:0] mesh_1_6_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177098.4]
  wire  mesh_1_6_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177098.4]
  wire [4:0] mesh_1_6_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177098.4]
  wire [7:0] mesh_1_6_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177098.4]
  wire [18:0] mesh_1_6_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177098.4]
  wire [18:0] mesh_1_6_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177098.4]
  wire  mesh_1_6_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177098.4]
  wire [4:0] mesh_1_6_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177098.4]
  wire  mesh_1_6_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177098.4]
  wire  mesh_1_6_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177098.4]
  wire  mesh_1_7_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177101.4]
  wire [7:0] mesh_1_7_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177101.4]
  wire [18:0] mesh_1_7_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177101.4]
  wire [18:0] mesh_1_7_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177101.4]
  wire  mesh_1_7_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177101.4]
  wire [4:0] mesh_1_7_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177101.4]
  wire [7:0] mesh_1_7_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177101.4]
  wire [18:0] mesh_1_7_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177101.4]
  wire [18:0] mesh_1_7_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177101.4]
  wire  mesh_1_7_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177101.4]
  wire [4:0] mesh_1_7_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177101.4]
  wire  mesh_1_7_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177101.4]
  wire  mesh_1_7_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177101.4]
  wire  mesh_2_0_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177104.4]
  wire [7:0] mesh_2_0_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177104.4]
  wire [18:0] mesh_2_0_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177104.4]
  wire [18:0] mesh_2_0_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177104.4]
  wire  mesh_2_0_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177104.4]
  wire [4:0] mesh_2_0_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177104.4]
  wire [7:0] mesh_2_0_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177104.4]
  wire [18:0] mesh_2_0_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177104.4]
  wire [18:0] mesh_2_0_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177104.4]
  wire  mesh_2_0_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177104.4]
  wire [4:0] mesh_2_0_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177104.4]
  wire  mesh_2_0_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177104.4]
  wire  mesh_2_0_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177104.4]
  wire  mesh_2_1_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177107.4]
  wire [7:0] mesh_2_1_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177107.4]
  wire [18:0] mesh_2_1_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177107.4]
  wire [18:0] mesh_2_1_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177107.4]
  wire  mesh_2_1_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177107.4]
  wire [4:0] mesh_2_1_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177107.4]
  wire [7:0] mesh_2_1_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177107.4]
  wire [18:0] mesh_2_1_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177107.4]
  wire [18:0] mesh_2_1_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177107.4]
  wire  mesh_2_1_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177107.4]
  wire [4:0] mesh_2_1_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177107.4]
  wire  mesh_2_1_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177107.4]
  wire  mesh_2_1_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177107.4]
  wire  mesh_2_2_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177110.4]
  wire [7:0] mesh_2_2_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177110.4]
  wire [18:0] mesh_2_2_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177110.4]
  wire [18:0] mesh_2_2_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177110.4]
  wire  mesh_2_2_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177110.4]
  wire [4:0] mesh_2_2_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177110.4]
  wire [7:0] mesh_2_2_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177110.4]
  wire [18:0] mesh_2_2_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177110.4]
  wire [18:0] mesh_2_2_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177110.4]
  wire  mesh_2_2_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177110.4]
  wire [4:0] mesh_2_2_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177110.4]
  wire  mesh_2_2_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177110.4]
  wire  mesh_2_2_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177110.4]
  wire  mesh_2_3_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177113.4]
  wire [7:0] mesh_2_3_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177113.4]
  wire [18:0] mesh_2_3_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177113.4]
  wire [18:0] mesh_2_3_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177113.4]
  wire  mesh_2_3_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177113.4]
  wire [4:0] mesh_2_3_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177113.4]
  wire [7:0] mesh_2_3_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177113.4]
  wire [18:0] mesh_2_3_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177113.4]
  wire [18:0] mesh_2_3_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177113.4]
  wire  mesh_2_3_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177113.4]
  wire [4:0] mesh_2_3_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177113.4]
  wire  mesh_2_3_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177113.4]
  wire  mesh_2_3_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177113.4]
  wire  mesh_2_4_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177116.4]
  wire [7:0] mesh_2_4_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177116.4]
  wire [18:0] mesh_2_4_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177116.4]
  wire [18:0] mesh_2_4_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177116.4]
  wire  mesh_2_4_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177116.4]
  wire [4:0] mesh_2_4_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177116.4]
  wire [7:0] mesh_2_4_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177116.4]
  wire [18:0] mesh_2_4_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177116.4]
  wire [18:0] mesh_2_4_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177116.4]
  wire  mesh_2_4_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177116.4]
  wire [4:0] mesh_2_4_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177116.4]
  wire  mesh_2_4_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177116.4]
  wire  mesh_2_4_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177116.4]
  wire  mesh_2_5_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177119.4]
  wire [7:0] mesh_2_5_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177119.4]
  wire [18:0] mesh_2_5_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177119.4]
  wire [18:0] mesh_2_5_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177119.4]
  wire  mesh_2_5_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177119.4]
  wire [4:0] mesh_2_5_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177119.4]
  wire [7:0] mesh_2_5_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177119.4]
  wire [18:0] mesh_2_5_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177119.4]
  wire [18:0] mesh_2_5_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177119.4]
  wire  mesh_2_5_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177119.4]
  wire [4:0] mesh_2_5_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177119.4]
  wire  mesh_2_5_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177119.4]
  wire  mesh_2_5_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177119.4]
  wire  mesh_2_6_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177122.4]
  wire [7:0] mesh_2_6_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177122.4]
  wire [18:0] mesh_2_6_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177122.4]
  wire [18:0] mesh_2_6_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177122.4]
  wire  mesh_2_6_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177122.4]
  wire [4:0] mesh_2_6_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177122.4]
  wire [7:0] mesh_2_6_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177122.4]
  wire [18:0] mesh_2_6_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177122.4]
  wire [18:0] mesh_2_6_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177122.4]
  wire  mesh_2_6_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177122.4]
  wire [4:0] mesh_2_6_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177122.4]
  wire  mesh_2_6_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177122.4]
  wire  mesh_2_6_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177122.4]
  wire  mesh_2_7_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177125.4]
  wire [7:0] mesh_2_7_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177125.4]
  wire [18:0] mesh_2_7_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177125.4]
  wire [18:0] mesh_2_7_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177125.4]
  wire  mesh_2_7_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177125.4]
  wire [4:0] mesh_2_7_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177125.4]
  wire [7:0] mesh_2_7_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177125.4]
  wire [18:0] mesh_2_7_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177125.4]
  wire [18:0] mesh_2_7_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177125.4]
  wire  mesh_2_7_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177125.4]
  wire [4:0] mesh_2_7_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177125.4]
  wire  mesh_2_7_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177125.4]
  wire  mesh_2_7_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177125.4]
  wire  mesh_3_0_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177128.4]
  wire [7:0] mesh_3_0_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177128.4]
  wire [18:0] mesh_3_0_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177128.4]
  wire [18:0] mesh_3_0_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177128.4]
  wire  mesh_3_0_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177128.4]
  wire [4:0] mesh_3_0_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177128.4]
  wire [7:0] mesh_3_0_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177128.4]
  wire [18:0] mesh_3_0_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177128.4]
  wire [18:0] mesh_3_0_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177128.4]
  wire  mesh_3_0_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177128.4]
  wire [4:0] mesh_3_0_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177128.4]
  wire  mesh_3_0_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177128.4]
  wire  mesh_3_0_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177128.4]
  wire  mesh_3_1_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177131.4]
  wire [7:0] mesh_3_1_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177131.4]
  wire [18:0] mesh_3_1_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177131.4]
  wire [18:0] mesh_3_1_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177131.4]
  wire  mesh_3_1_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177131.4]
  wire [4:0] mesh_3_1_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177131.4]
  wire [7:0] mesh_3_1_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177131.4]
  wire [18:0] mesh_3_1_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177131.4]
  wire [18:0] mesh_3_1_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177131.4]
  wire  mesh_3_1_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177131.4]
  wire [4:0] mesh_3_1_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177131.4]
  wire  mesh_3_1_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177131.4]
  wire  mesh_3_1_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177131.4]
  wire  mesh_3_2_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177134.4]
  wire [7:0] mesh_3_2_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177134.4]
  wire [18:0] mesh_3_2_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177134.4]
  wire [18:0] mesh_3_2_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177134.4]
  wire  mesh_3_2_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177134.4]
  wire [4:0] mesh_3_2_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177134.4]
  wire [7:0] mesh_3_2_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177134.4]
  wire [18:0] mesh_3_2_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177134.4]
  wire [18:0] mesh_3_2_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177134.4]
  wire  mesh_3_2_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177134.4]
  wire [4:0] mesh_3_2_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177134.4]
  wire  mesh_3_2_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177134.4]
  wire  mesh_3_2_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177134.4]
  wire  mesh_3_3_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177137.4]
  wire [7:0] mesh_3_3_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177137.4]
  wire [18:0] mesh_3_3_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177137.4]
  wire [18:0] mesh_3_3_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177137.4]
  wire  mesh_3_3_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177137.4]
  wire [4:0] mesh_3_3_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177137.4]
  wire [7:0] mesh_3_3_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177137.4]
  wire [18:0] mesh_3_3_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177137.4]
  wire [18:0] mesh_3_3_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177137.4]
  wire  mesh_3_3_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177137.4]
  wire [4:0] mesh_3_3_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177137.4]
  wire  mesh_3_3_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177137.4]
  wire  mesh_3_3_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177137.4]
  wire  mesh_3_4_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177140.4]
  wire [7:0] mesh_3_4_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177140.4]
  wire [18:0] mesh_3_4_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177140.4]
  wire [18:0] mesh_3_4_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177140.4]
  wire  mesh_3_4_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177140.4]
  wire [4:0] mesh_3_4_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177140.4]
  wire [7:0] mesh_3_4_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177140.4]
  wire [18:0] mesh_3_4_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177140.4]
  wire [18:0] mesh_3_4_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177140.4]
  wire  mesh_3_4_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177140.4]
  wire [4:0] mesh_3_4_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177140.4]
  wire  mesh_3_4_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177140.4]
  wire  mesh_3_4_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177140.4]
  wire  mesh_3_5_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177143.4]
  wire [7:0] mesh_3_5_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177143.4]
  wire [18:0] mesh_3_5_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177143.4]
  wire [18:0] mesh_3_5_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177143.4]
  wire  mesh_3_5_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177143.4]
  wire [4:0] mesh_3_5_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177143.4]
  wire [7:0] mesh_3_5_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177143.4]
  wire [18:0] mesh_3_5_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177143.4]
  wire [18:0] mesh_3_5_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177143.4]
  wire  mesh_3_5_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177143.4]
  wire [4:0] mesh_3_5_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177143.4]
  wire  mesh_3_5_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177143.4]
  wire  mesh_3_5_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177143.4]
  wire  mesh_3_6_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177146.4]
  wire [7:0] mesh_3_6_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177146.4]
  wire [18:0] mesh_3_6_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177146.4]
  wire [18:0] mesh_3_6_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177146.4]
  wire  mesh_3_6_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177146.4]
  wire [4:0] mesh_3_6_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177146.4]
  wire [7:0] mesh_3_6_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177146.4]
  wire [18:0] mesh_3_6_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177146.4]
  wire [18:0] mesh_3_6_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177146.4]
  wire  mesh_3_6_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177146.4]
  wire [4:0] mesh_3_6_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177146.4]
  wire  mesh_3_6_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177146.4]
  wire  mesh_3_6_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177146.4]
  wire  mesh_3_7_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177149.4]
  wire [7:0] mesh_3_7_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177149.4]
  wire [18:0] mesh_3_7_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177149.4]
  wire [18:0] mesh_3_7_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177149.4]
  wire  mesh_3_7_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177149.4]
  wire [4:0] mesh_3_7_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177149.4]
  wire [7:0] mesh_3_7_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177149.4]
  wire [18:0] mesh_3_7_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177149.4]
  wire [18:0] mesh_3_7_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177149.4]
  wire  mesh_3_7_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177149.4]
  wire [4:0] mesh_3_7_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177149.4]
  wire  mesh_3_7_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177149.4]
  wire  mesh_3_7_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177149.4]
  wire  mesh_4_0_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177152.4]
  wire [7:0] mesh_4_0_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177152.4]
  wire [18:0] mesh_4_0_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177152.4]
  wire [18:0] mesh_4_0_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177152.4]
  wire  mesh_4_0_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177152.4]
  wire [4:0] mesh_4_0_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177152.4]
  wire [7:0] mesh_4_0_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177152.4]
  wire [18:0] mesh_4_0_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177152.4]
  wire [18:0] mesh_4_0_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177152.4]
  wire  mesh_4_0_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177152.4]
  wire [4:0] mesh_4_0_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177152.4]
  wire  mesh_4_0_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177152.4]
  wire  mesh_4_0_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177152.4]
  wire  mesh_4_1_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177155.4]
  wire [7:0] mesh_4_1_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177155.4]
  wire [18:0] mesh_4_1_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177155.4]
  wire [18:0] mesh_4_1_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177155.4]
  wire  mesh_4_1_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177155.4]
  wire [4:0] mesh_4_1_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177155.4]
  wire [7:0] mesh_4_1_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177155.4]
  wire [18:0] mesh_4_1_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177155.4]
  wire [18:0] mesh_4_1_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177155.4]
  wire  mesh_4_1_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177155.4]
  wire [4:0] mesh_4_1_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177155.4]
  wire  mesh_4_1_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177155.4]
  wire  mesh_4_1_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177155.4]
  wire  mesh_4_2_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177158.4]
  wire [7:0] mesh_4_2_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177158.4]
  wire [18:0] mesh_4_2_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177158.4]
  wire [18:0] mesh_4_2_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177158.4]
  wire  mesh_4_2_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177158.4]
  wire [4:0] mesh_4_2_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177158.4]
  wire [7:0] mesh_4_2_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177158.4]
  wire [18:0] mesh_4_2_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177158.4]
  wire [18:0] mesh_4_2_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177158.4]
  wire  mesh_4_2_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177158.4]
  wire [4:0] mesh_4_2_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177158.4]
  wire  mesh_4_2_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177158.4]
  wire  mesh_4_2_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177158.4]
  wire  mesh_4_3_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177161.4]
  wire [7:0] mesh_4_3_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177161.4]
  wire [18:0] mesh_4_3_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177161.4]
  wire [18:0] mesh_4_3_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177161.4]
  wire  mesh_4_3_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177161.4]
  wire [4:0] mesh_4_3_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177161.4]
  wire [7:0] mesh_4_3_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177161.4]
  wire [18:0] mesh_4_3_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177161.4]
  wire [18:0] mesh_4_3_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177161.4]
  wire  mesh_4_3_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177161.4]
  wire [4:0] mesh_4_3_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177161.4]
  wire  mesh_4_3_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177161.4]
  wire  mesh_4_3_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177161.4]
  wire  mesh_4_4_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177164.4]
  wire [7:0] mesh_4_4_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177164.4]
  wire [18:0] mesh_4_4_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177164.4]
  wire [18:0] mesh_4_4_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177164.4]
  wire  mesh_4_4_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177164.4]
  wire [4:0] mesh_4_4_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177164.4]
  wire [7:0] mesh_4_4_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177164.4]
  wire [18:0] mesh_4_4_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177164.4]
  wire [18:0] mesh_4_4_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177164.4]
  wire  mesh_4_4_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177164.4]
  wire [4:0] mesh_4_4_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177164.4]
  wire  mesh_4_4_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177164.4]
  wire  mesh_4_4_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177164.4]
  wire  mesh_4_5_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177167.4]
  wire [7:0] mesh_4_5_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177167.4]
  wire [18:0] mesh_4_5_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177167.4]
  wire [18:0] mesh_4_5_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177167.4]
  wire  mesh_4_5_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177167.4]
  wire [4:0] mesh_4_5_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177167.4]
  wire [7:0] mesh_4_5_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177167.4]
  wire [18:0] mesh_4_5_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177167.4]
  wire [18:0] mesh_4_5_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177167.4]
  wire  mesh_4_5_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177167.4]
  wire [4:0] mesh_4_5_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177167.4]
  wire  mesh_4_5_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177167.4]
  wire  mesh_4_5_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177167.4]
  wire  mesh_4_6_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177170.4]
  wire [7:0] mesh_4_6_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177170.4]
  wire [18:0] mesh_4_6_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177170.4]
  wire [18:0] mesh_4_6_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177170.4]
  wire  mesh_4_6_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177170.4]
  wire [4:0] mesh_4_6_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177170.4]
  wire [7:0] mesh_4_6_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177170.4]
  wire [18:0] mesh_4_6_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177170.4]
  wire [18:0] mesh_4_6_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177170.4]
  wire  mesh_4_6_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177170.4]
  wire [4:0] mesh_4_6_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177170.4]
  wire  mesh_4_6_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177170.4]
  wire  mesh_4_6_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177170.4]
  wire  mesh_4_7_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177173.4]
  wire [7:0] mesh_4_7_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177173.4]
  wire [18:0] mesh_4_7_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177173.4]
  wire [18:0] mesh_4_7_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177173.4]
  wire  mesh_4_7_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177173.4]
  wire [4:0] mesh_4_7_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177173.4]
  wire [7:0] mesh_4_7_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177173.4]
  wire [18:0] mesh_4_7_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177173.4]
  wire [18:0] mesh_4_7_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177173.4]
  wire  mesh_4_7_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177173.4]
  wire [4:0] mesh_4_7_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177173.4]
  wire  mesh_4_7_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177173.4]
  wire  mesh_4_7_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177173.4]
  wire  mesh_5_0_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177176.4]
  wire [7:0] mesh_5_0_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177176.4]
  wire [18:0] mesh_5_0_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177176.4]
  wire [18:0] mesh_5_0_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177176.4]
  wire  mesh_5_0_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177176.4]
  wire [4:0] mesh_5_0_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177176.4]
  wire [7:0] mesh_5_0_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177176.4]
  wire [18:0] mesh_5_0_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177176.4]
  wire [18:0] mesh_5_0_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177176.4]
  wire  mesh_5_0_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177176.4]
  wire [4:0] mesh_5_0_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177176.4]
  wire  mesh_5_0_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177176.4]
  wire  mesh_5_0_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177176.4]
  wire  mesh_5_1_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177179.4]
  wire [7:0] mesh_5_1_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177179.4]
  wire [18:0] mesh_5_1_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177179.4]
  wire [18:0] mesh_5_1_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177179.4]
  wire  mesh_5_1_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177179.4]
  wire [4:0] mesh_5_1_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177179.4]
  wire [7:0] mesh_5_1_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177179.4]
  wire [18:0] mesh_5_1_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177179.4]
  wire [18:0] mesh_5_1_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177179.4]
  wire  mesh_5_1_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177179.4]
  wire [4:0] mesh_5_1_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177179.4]
  wire  mesh_5_1_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177179.4]
  wire  mesh_5_1_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177179.4]
  wire  mesh_5_2_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177182.4]
  wire [7:0] mesh_5_2_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177182.4]
  wire [18:0] mesh_5_2_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177182.4]
  wire [18:0] mesh_5_2_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177182.4]
  wire  mesh_5_2_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177182.4]
  wire [4:0] mesh_5_2_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177182.4]
  wire [7:0] mesh_5_2_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177182.4]
  wire [18:0] mesh_5_2_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177182.4]
  wire [18:0] mesh_5_2_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177182.4]
  wire  mesh_5_2_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177182.4]
  wire [4:0] mesh_5_2_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177182.4]
  wire  mesh_5_2_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177182.4]
  wire  mesh_5_2_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177182.4]
  wire  mesh_5_3_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177185.4]
  wire [7:0] mesh_5_3_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177185.4]
  wire [18:0] mesh_5_3_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177185.4]
  wire [18:0] mesh_5_3_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177185.4]
  wire  mesh_5_3_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177185.4]
  wire [4:0] mesh_5_3_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177185.4]
  wire [7:0] mesh_5_3_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177185.4]
  wire [18:0] mesh_5_3_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177185.4]
  wire [18:0] mesh_5_3_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177185.4]
  wire  mesh_5_3_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177185.4]
  wire [4:0] mesh_5_3_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177185.4]
  wire  mesh_5_3_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177185.4]
  wire  mesh_5_3_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177185.4]
  wire  mesh_5_4_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177188.4]
  wire [7:0] mesh_5_4_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177188.4]
  wire [18:0] mesh_5_4_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177188.4]
  wire [18:0] mesh_5_4_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177188.4]
  wire  mesh_5_4_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177188.4]
  wire [4:0] mesh_5_4_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177188.4]
  wire [7:0] mesh_5_4_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177188.4]
  wire [18:0] mesh_5_4_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177188.4]
  wire [18:0] mesh_5_4_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177188.4]
  wire  mesh_5_4_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177188.4]
  wire [4:0] mesh_5_4_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177188.4]
  wire  mesh_5_4_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177188.4]
  wire  mesh_5_4_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177188.4]
  wire  mesh_5_5_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177191.4]
  wire [7:0] mesh_5_5_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177191.4]
  wire [18:0] mesh_5_5_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177191.4]
  wire [18:0] mesh_5_5_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177191.4]
  wire  mesh_5_5_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177191.4]
  wire [4:0] mesh_5_5_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177191.4]
  wire [7:0] mesh_5_5_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177191.4]
  wire [18:0] mesh_5_5_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177191.4]
  wire [18:0] mesh_5_5_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177191.4]
  wire  mesh_5_5_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177191.4]
  wire [4:0] mesh_5_5_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177191.4]
  wire  mesh_5_5_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177191.4]
  wire  mesh_5_5_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177191.4]
  wire  mesh_5_6_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177194.4]
  wire [7:0] mesh_5_6_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177194.4]
  wire [18:0] mesh_5_6_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177194.4]
  wire [18:0] mesh_5_6_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177194.4]
  wire  mesh_5_6_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177194.4]
  wire [4:0] mesh_5_6_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177194.4]
  wire [7:0] mesh_5_6_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177194.4]
  wire [18:0] mesh_5_6_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177194.4]
  wire [18:0] mesh_5_6_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177194.4]
  wire  mesh_5_6_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177194.4]
  wire [4:0] mesh_5_6_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177194.4]
  wire  mesh_5_6_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177194.4]
  wire  mesh_5_6_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177194.4]
  wire  mesh_5_7_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177197.4]
  wire [7:0] mesh_5_7_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177197.4]
  wire [18:0] mesh_5_7_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177197.4]
  wire [18:0] mesh_5_7_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177197.4]
  wire  mesh_5_7_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177197.4]
  wire [4:0] mesh_5_7_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177197.4]
  wire [7:0] mesh_5_7_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177197.4]
  wire [18:0] mesh_5_7_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177197.4]
  wire [18:0] mesh_5_7_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177197.4]
  wire  mesh_5_7_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177197.4]
  wire [4:0] mesh_5_7_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177197.4]
  wire  mesh_5_7_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177197.4]
  wire  mesh_5_7_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177197.4]
  wire  mesh_6_0_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177200.4]
  wire [7:0] mesh_6_0_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177200.4]
  wire [18:0] mesh_6_0_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177200.4]
  wire [18:0] mesh_6_0_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177200.4]
  wire  mesh_6_0_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177200.4]
  wire [4:0] mesh_6_0_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177200.4]
  wire [7:0] mesh_6_0_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177200.4]
  wire [18:0] mesh_6_0_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177200.4]
  wire [18:0] mesh_6_0_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177200.4]
  wire  mesh_6_0_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177200.4]
  wire [4:0] mesh_6_0_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177200.4]
  wire  mesh_6_0_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177200.4]
  wire  mesh_6_0_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177200.4]
  wire  mesh_6_1_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177203.4]
  wire [7:0] mesh_6_1_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177203.4]
  wire [18:0] mesh_6_1_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177203.4]
  wire [18:0] mesh_6_1_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177203.4]
  wire  mesh_6_1_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177203.4]
  wire [4:0] mesh_6_1_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177203.4]
  wire [7:0] mesh_6_1_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177203.4]
  wire [18:0] mesh_6_1_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177203.4]
  wire [18:0] mesh_6_1_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177203.4]
  wire  mesh_6_1_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177203.4]
  wire [4:0] mesh_6_1_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177203.4]
  wire  mesh_6_1_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177203.4]
  wire  mesh_6_1_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177203.4]
  wire  mesh_6_2_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177206.4]
  wire [7:0] mesh_6_2_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177206.4]
  wire [18:0] mesh_6_2_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177206.4]
  wire [18:0] mesh_6_2_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177206.4]
  wire  mesh_6_2_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177206.4]
  wire [4:0] mesh_6_2_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177206.4]
  wire [7:0] mesh_6_2_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177206.4]
  wire [18:0] mesh_6_2_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177206.4]
  wire [18:0] mesh_6_2_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177206.4]
  wire  mesh_6_2_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177206.4]
  wire [4:0] mesh_6_2_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177206.4]
  wire  mesh_6_2_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177206.4]
  wire  mesh_6_2_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177206.4]
  wire  mesh_6_3_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177209.4]
  wire [7:0] mesh_6_3_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177209.4]
  wire [18:0] mesh_6_3_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177209.4]
  wire [18:0] mesh_6_3_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177209.4]
  wire  mesh_6_3_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177209.4]
  wire [4:0] mesh_6_3_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177209.4]
  wire [7:0] mesh_6_3_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177209.4]
  wire [18:0] mesh_6_3_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177209.4]
  wire [18:0] mesh_6_3_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177209.4]
  wire  mesh_6_3_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177209.4]
  wire [4:0] mesh_6_3_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177209.4]
  wire  mesh_6_3_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177209.4]
  wire  mesh_6_3_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177209.4]
  wire  mesh_6_4_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177212.4]
  wire [7:0] mesh_6_4_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177212.4]
  wire [18:0] mesh_6_4_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177212.4]
  wire [18:0] mesh_6_4_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177212.4]
  wire  mesh_6_4_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177212.4]
  wire [4:0] mesh_6_4_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177212.4]
  wire [7:0] mesh_6_4_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177212.4]
  wire [18:0] mesh_6_4_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177212.4]
  wire [18:0] mesh_6_4_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177212.4]
  wire  mesh_6_4_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177212.4]
  wire [4:0] mesh_6_4_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177212.4]
  wire  mesh_6_4_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177212.4]
  wire  mesh_6_4_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177212.4]
  wire  mesh_6_5_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177215.4]
  wire [7:0] mesh_6_5_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177215.4]
  wire [18:0] mesh_6_5_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177215.4]
  wire [18:0] mesh_6_5_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177215.4]
  wire  mesh_6_5_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177215.4]
  wire [4:0] mesh_6_5_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177215.4]
  wire [7:0] mesh_6_5_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177215.4]
  wire [18:0] mesh_6_5_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177215.4]
  wire [18:0] mesh_6_5_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177215.4]
  wire  mesh_6_5_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177215.4]
  wire [4:0] mesh_6_5_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177215.4]
  wire  mesh_6_5_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177215.4]
  wire  mesh_6_5_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177215.4]
  wire  mesh_6_6_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177218.4]
  wire [7:0] mesh_6_6_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177218.4]
  wire [18:0] mesh_6_6_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177218.4]
  wire [18:0] mesh_6_6_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177218.4]
  wire  mesh_6_6_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177218.4]
  wire [4:0] mesh_6_6_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177218.4]
  wire [7:0] mesh_6_6_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177218.4]
  wire [18:0] mesh_6_6_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177218.4]
  wire [18:0] mesh_6_6_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177218.4]
  wire  mesh_6_6_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177218.4]
  wire [4:0] mesh_6_6_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177218.4]
  wire  mesh_6_6_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177218.4]
  wire  mesh_6_6_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177218.4]
  wire  mesh_6_7_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177221.4]
  wire [7:0] mesh_6_7_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177221.4]
  wire [18:0] mesh_6_7_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177221.4]
  wire [18:0] mesh_6_7_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177221.4]
  wire  mesh_6_7_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177221.4]
  wire [4:0] mesh_6_7_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177221.4]
  wire [7:0] mesh_6_7_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177221.4]
  wire [18:0] mesh_6_7_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177221.4]
  wire [18:0] mesh_6_7_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177221.4]
  wire  mesh_6_7_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177221.4]
  wire [4:0] mesh_6_7_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177221.4]
  wire  mesh_6_7_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177221.4]
  wire  mesh_6_7_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177221.4]
  wire  mesh_7_0_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177224.4]
  wire [7:0] mesh_7_0_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177224.4]
  wire [18:0] mesh_7_0_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177224.4]
  wire [18:0] mesh_7_0_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177224.4]
  wire  mesh_7_0_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177224.4]
  wire [4:0] mesh_7_0_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177224.4]
  wire [7:0] mesh_7_0_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177224.4]
  wire [18:0] mesh_7_0_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177224.4]
  wire [18:0] mesh_7_0_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177224.4]
  wire  mesh_7_0_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177224.4]
  wire [4:0] mesh_7_0_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177224.4]
  wire  mesh_7_0_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177224.4]
  wire  mesh_7_0_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177224.4]
  wire  mesh_7_1_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177227.4]
  wire [7:0] mesh_7_1_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177227.4]
  wire [18:0] mesh_7_1_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177227.4]
  wire [18:0] mesh_7_1_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177227.4]
  wire  mesh_7_1_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177227.4]
  wire [4:0] mesh_7_1_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177227.4]
  wire [7:0] mesh_7_1_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177227.4]
  wire [18:0] mesh_7_1_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177227.4]
  wire [18:0] mesh_7_1_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177227.4]
  wire  mesh_7_1_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177227.4]
  wire [4:0] mesh_7_1_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177227.4]
  wire  mesh_7_1_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177227.4]
  wire  mesh_7_1_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177227.4]
  wire  mesh_7_2_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177230.4]
  wire [7:0] mesh_7_2_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177230.4]
  wire [18:0] mesh_7_2_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177230.4]
  wire [18:0] mesh_7_2_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177230.4]
  wire  mesh_7_2_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177230.4]
  wire [4:0] mesh_7_2_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177230.4]
  wire [7:0] mesh_7_2_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177230.4]
  wire [18:0] mesh_7_2_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177230.4]
  wire [18:0] mesh_7_2_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177230.4]
  wire  mesh_7_2_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177230.4]
  wire [4:0] mesh_7_2_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177230.4]
  wire  mesh_7_2_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177230.4]
  wire  mesh_7_2_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177230.4]
  wire  mesh_7_3_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177233.4]
  wire [7:0] mesh_7_3_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177233.4]
  wire [18:0] mesh_7_3_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177233.4]
  wire [18:0] mesh_7_3_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177233.4]
  wire  mesh_7_3_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177233.4]
  wire [4:0] mesh_7_3_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177233.4]
  wire [7:0] mesh_7_3_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177233.4]
  wire [18:0] mesh_7_3_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177233.4]
  wire [18:0] mesh_7_3_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177233.4]
  wire  mesh_7_3_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177233.4]
  wire [4:0] mesh_7_3_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177233.4]
  wire  mesh_7_3_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177233.4]
  wire  mesh_7_3_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177233.4]
  wire  mesh_7_4_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177236.4]
  wire [7:0] mesh_7_4_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177236.4]
  wire [18:0] mesh_7_4_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177236.4]
  wire [18:0] mesh_7_4_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177236.4]
  wire  mesh_7_4_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177236.4]
  wire [4:0] mesh_7_4_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177236.4]
  wire [7:0] mesh_7_4_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177236.4]
  wire [18:0] mesh_7_4_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177236.4]
  wire [18:0] mesh_7_4_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177236.4]
  wire  mesh_7_4_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177236.4]
  wire [4:0] mesh_7_4_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177236.4]
  wire  mesh_7_4_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177236.4]
  wire  mesh_7_4_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177236.4]
  wire  mesh_7_5_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177239.4]
  wire [7:0] mesh_7_5_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177239.4]
  wire [18:0] mesh_7_5_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177239.4]
  wire [18:0] mesh_7_5_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177239.4]
  wire  mesh_7_5_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177239.4]
  wire [4:0] mesh_7_5_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177239.4]
  wire [7:0] mesh_7_5_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177239.4]
  wire [18:0] mesh_7_5_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177239.4]
  wire [18:0] mesh_7_5_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177239.4]
  wire  mesh_7_5_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177239.4]
  wire [4:0] mesh_7_5_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177239.4]
  wire  mesh_7_5_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177239.4]
  wire  mesh_7_5_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177239.4]
  wire  mesh_7_6_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177242.4]
  wire [7:0] mesh_7_6_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177242.4]
  wire [18:0] mesh_7_6_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177242.4]
  wire [18:0] mesh_7_6_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177242.4]
  wire  mesh_7_6_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177242.4]
  wire [4:0] mesh_7_6_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177242.4]
  wire [7:0] mesh_7_6_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177242.4]
  wire [18:0] mesh_7_6_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177242.4]
  wire [18:0] mesh_7_6_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177242.4]
  wire  mesh_7_6_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177242.4]
  wire [4:0] mesh_7_6_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177242.4]
  wire  mesh_7_6_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177242.4]
  wire  mesh_7_6_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177242.4]
  wire  mesh_7_7_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177245.4]
  wire [7:0] mesh_7_7_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177245.4]
  wire [18:0] mesh_7_7_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177245.4]
  wire [18:0] mesh_7_7_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177245.4]
  wire  mesh_7_7_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177245.4]
  wire [4:0] mesh_7_7_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177245.4]
  wire [7:0] mesh_7_7_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177245.4]
  wire [18:0] mesh_7_7_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177245.4]
  wire [18:0] mesh_7_7_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177245.4]
  wire  mesh_7_7_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177245.4]
  wire [4:0] mesh_7_7_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177245.4]
  wire  mesh_7_7_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177245.4]
  wire  mesh_7_7_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177245.4]
  reg [7:0] _T_0; // @[Mesh.scala 40:29:example.TestHarness.GemminiSocTest1RocketConfig.fir@177248.4]
  reg [31:0] _RAND_0;
  reg [7:0] _T_1_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177250.4]
  reg [31:0] _RAND_1;
  reg [7:0] _T_2_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177253.4]
  reg [31:0] _RAND_2;
  reg [7:0] _T_3_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177256.4]
  reg [31:0] _RAND_3;
  reg [7:0] _T_4_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177259.4]
  reg [31:0] _RAND_4;
  reg [7:0] _T_5_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177262.4]
  reg [31:0] _RAND_5;
  reg [7:0] _T_6_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177265.4]
  reg [31:0] _RAND_6;
  reg [7:0] _T_7_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177268.4]
  reg [31:0] _RAND_7;
  reg [7:0] _T_8_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177271.4]
  reg [31:0] _RAND_8;
  reg [7:0] _T_9_0; // @[Mesh.scala 40:29:example.TestHarness.GemminiSocTest1RocketConfig.fir@177274.4]
  reg [31:0] _RAND_9;
  reg [7:0] _T_10_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177276.4]
  reg [31:0] _RAND_10;
  reg [7:0] _T_11_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177279.4]
  reg [31:0] _RAND_11;
  reg [7:0] _T_12_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177282.4]
  reg [31:0] _RAND_12;
  reg [7:0] _T_13_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177285.4]
  reg [31:0] _RAND_13;
  reg [7:0] _T_14_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177288.4]
  reg [31:0] _RAND_14;
  reg [7:0] _T_15_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177291.4]
  reg [31:0] _RAND_15;
  reg [7:0] _T_16_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177294.4]
  reg [31:0] _RAND_16;
  reg [7:0] _T_17_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177297.4]
  reg [31:0] _RAND_17;
  reg [7:0] _T_18_0; // @[Mesh.scala 40:29:example.TestHarness.GemminiSocTest1RocketConfig.fir@177300.4]
  reg [31:0] _RAND_18;
  reg [7:0] _T_19_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177302.4]
  reg [31:0] _RAND_19;
  reg [7:0] _T_20_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177305.4]
  reg [31:0] _RAND_20;
  reg [7:0] _T_21_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177308.4]
  reg [31:0] _RAND_21;
  reg [7:0] _T_22_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177311.4]
  reg [31:0] _RAND_22;
  reg [7:0] _T_23_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177314.4]
  reg [31:0] _RAND_23;
  reg [7:0] _T_24_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177317.4]
  reg [31:0] _RAND_24;
  reg [7:0] _T_25_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177320.4]
  reg [31:0] _RAND_25;
  reg [7:0] _T_26_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177323.4]
  reg [31:0] _RAND_26;
  reg [7:0] _T_27_0; // @[Mesh.scala 40:29:example.TestHarness.GemminiSocTest1RocketConfig.fir@177326.4]
  reg [31:0] _RAND_27;
  reg [7:0] _T_28_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177328.4]
  reg [31:0] _RAND_28;
  reg [7:0] _T_29_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177331.4]
  reg [31:0] _RAND_29;
  reg [7:0] _T_30_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177334.4]
  reg [31:0] _RAND_30;
  reg [7:0] _T_31_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177337.4]
  reg [31:0] _RAND_31;
  reg [7:0] _T_32_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177340.4]
  reg [31:0] _RAND_32;
  reg [7:0] _T_33_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177343.4]
  reg [31:0] _RAND_33;
  reg [7:0] _T_34_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177346.4]
  reg [31:0] _RAND_34;
  reg [7:0] _T_35_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177349.4]
  reg [31:0] _RAND_35;
  reg [7:0] _T_36_0; // @[Mesh.scala 40:29:example.TestHarness.GemminiSocTest1RocketConfig.fir@177352.4]
  reg [31:0] _RAND_36;
  reg [7:0] _T_37_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177354.4]
  reg [31:0] _RAND_37;
  reg [7:0] _T_38_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177357.4]
  reg [31:0] _RAND_38;
  reg [7:0] _T_39_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177360.4]
  reg [31:0] _RAND_39;
  reg [7:0] _T_40_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177363.4]
  reg [31:0] _RAND_40;
  reg [7:0] _T_41_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177366.4]
  reg [31:0] _RAND_41;
  reg [7:0] _T_42_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177369.4]
  reg [31:0] _RAND_42;
  reg [7:0] _T_43_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177372.4]
  reg [31:0] _RAND_43;
  reg [7:0] _T_44_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177375.4]
  reg [31:0] _RAND_44;
  reg [7:0] _T_45_0; // @[Mesh.scala 40:29:example.TestHarness.GemminiSocTest1RocketConfig.fir@177378.4]
  reg [31:0] _RAND_45;
  reg [7:0] _T_46_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177380.4]
  reg [31:0] _RAND_46;
  reg [7:0] _T_47_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177383.4]
  reg [31:0] _RAND_47;
  reg [7:0] _T_48_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177386.4]
  reg [31:0] _RAND_48;
  reg [7:0] _T_49_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177389.4]
  reg [31:0] _RAND_49;
  reg [7:0] _T_50_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177392.4]
  reg [31:0] _RAND_50;
  reg [7:0] _T_51_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177395.4]
  reg [31:0] _RAND_51;
  reg [7:0] _T_52_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177398.4]
  reg [31:0] _RAND_52;
  reg [7:0] _T_53_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177401.4]
  reg [31:0] _RAND_53;
  reg [7:0] _T_54_0; // @[Mesh.scala 40:29:example.TestHarness.GemminiSocTest1RocketConfig.fir@177404.4]
  reg [31:0] _RAND_54;
  reg [7:0] _T_55_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177406.4]
  reg [31:0] _RAND_55;
  reg [7:0] _T_56_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177409.4]
  reg [31:0] _RAND_56;
  reg [7:0] _T_57_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177412.4]
  reg [31:0] _RAND_57;
  reg [7:0] _T_58_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177415.4]
  reg [31:0] _RAND_58;
  reg [7:0] _T_59_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177418.4]
  reg [31:0] _RAND_59;
  reg [7:0] _T_60_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177421.4]
  reg [31:0] _RAND_60;
  reg [7:0] _T_61_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177424.4]
  reg [31:0] _RAND_61;
  reg [7:0] _T_62_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177427.4]
  reg [31:0] _RAND_62;
  reg [7:0] _T_63_0; // @[Mesh.scala 40:29:example.TestHarness.GemminiSocTest1RocketConfig.fir@177430.4]
  reg [31:0] _RAND_63;
  reg [7:0] _T_64_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177432.4]
  reg [31:0] _RAND_64;
  reg [7:0] _T_65_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177435.4]
  reg [31:0] _RAND_65;
  reg [7:0] _T_66_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177438.4]
  reg [31:0] _RAND_66;
  reg [7:0] _T_67_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177441.4]
  reg [31:0] _RAND_67;
  reg [7:0] _T_68_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177444.4]
  reg [31:0] _RAND_68;
  reg [7:0] _T_69_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177447.4]
  reg [31:0] _RAND_69;
  reg [7:0] _T_70_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177450.4]
  reg [31:0] _RAND_70;
  reg [7:0] _T_71_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig.fir@177453.4]
  reg [31:0] _RAND_71;
  reg [7:0] _T_72_0; // @[Mesh.scala 48:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@177456.4]
  reg [31:0] _RAND_72;
  reg  _T_73_0; // @[Mesh.scala 48:52:example.TestHarness.GemminiSocTest1RocketConfig.fir@177458.4]
  reg [31:0] _RAND_73;
  reg [7:0] _T_74_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177460.4]
  reg [31:0] _RAND_74;
  reg [18:0] _T_75_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177465.4]
  reg [31:0] _RAND_75;
  reg [18:0] _T_76_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177470.4]
  reg [31:0] _RAND_76;
  reg [18:0] _T_77_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177475.4]
  reg [31:0] _RAND_77;
  reg [18:0] _T_78_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177480.4]
  reg [31:0] _RAND_78;
  reg [18:0] _T_79_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177485.4]
  reg [31:0] _RAND_79;
  reg [18:0] _T_80_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177490.4]
  reg [31:0] _RAND_80;
  reg [18:0] _T_81_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177495.4]
  reg [31:0] _RAND_81;
  reg [7:0] _T_82_0; // @[Mesh.scala 48:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@177500.4]
  reg [31:0] _RAND_82;
  reg  _T_83_0; // @[Mesh.scala 48:52:example.TestHarness.GemminiSocTest1RocketConfig.fir@177502.4]
  reg [31:0] _RAND_83;
  reg [7:0] _T_84_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177504.4]
  reg [31:0] _RAND_84;
  reg [18:0] _T_85_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177509.4]
  reg [31:0] _RAND_85;
  reg [18:0] _T_86_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177514.4]
  reg [31:0] _RAND_86;
  reg [18:0] _T_87_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177519.4]
  reg [31:0] _RAND_87;
  reg [18:0] _T_88_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177524.4]
  reg [31:0] _RAND_88;
  reg [18:0] _T_89_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177529.4]
  reg [31:0] _RAND_89;
  reg [18:0] _T_90_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177534.4]
  reg [31:0] _RAND_90;
  reg [18:0] _T_91_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177539.4]
  reg [31:0] _RAND_91;
  reg [7:0] _T_92_0; // @[Mesh.scala 48:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@177544.4]
  reg [31:0] _RAND_92;
  reg  _T_93_0; // @[Mesh.scala 48:52:example.TestHarness.GemminiSocTest1RocketConfig.fir@177546.4]
  reg [31:0] _RAND_93;
  reg [7:0] _T_94_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177548.4]
  reg [31:0] _RAND_94;
  reg [18:0] _T_95_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177553.4]
  reg [31:0] _RAND_95;
  reg [18:0] _T_96_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177558.4]
  reg [31:0] _RAND_96;
  reg [18:0] _T_97_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177563.4]
  reg [31:0] _RAND_97;
  reg [18:0] _T_98_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177568.4]
  reg [31:0] _RAND_98;
  reg [18:0] _T_99_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177573.4]
  reg [31:0] _RAND_99;
  reg [18:0] _T_100_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177578.4]
  reg [31:0] _RAND_100;
  reg [18:0] _T_101_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177583.4]
  reg [31:0] _RAND_101;
  reg [7:0] _T_102_0; // @[Mesh.scala 48:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@177588.4]
  reg [31:0] _RAND_102;
  reg  _T_103_0; // @[Mesh.scala 48:52:example.TestHarness.GemminiSocTest1RocketConfig.fir@177590.4]
  reg [31:0] _RAND_103;
  reg [7:0] _T_104_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177592.4]
  reg [31:0] _RAND_104;
  reg [18:0] _T_105_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177597.4]
  reg [31:0] _RAND_105;
  reg [18:0] _T_106_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177602.4]
  reg [31:0] _RAND_106;
  reg [18:0] _T_107_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177607.4]
  reg [31:0] _RAND_107;
  reg [18:0] _T_108_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177612.4]
  reg [31:0] _RAND_108;
  reg [18:0] _T_109_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177617.4]
  reg [31:0] _RAND_109;
  reg [18:0] _T_110_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177622.4]
  reg [31:0] _RAND_110;
  reg [18:0] _T_111_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177627.4]
  reg [31:0] _RAND_111;
  reg [7:0] _T_112_0; // @[Mesh.scala 48:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@177632.4]
  reg [31:0] _RAND_112;
  reg  _T_113_0; // @[Mesh.scala 48:52:example.TestHarness.GemminiSocTest1RocketConfig.fir@177634.4]
  reg [31:0] _RAND_113;
  reg [7:0] _T_114_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177636.4]
  reg [31:0] _RAND_114;
  reg [18:0] _T_115_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177641.4]
  reg [31:0] _RAND_115;
  reg [18:0] _T_116_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177646.4]
  reg [31:0] _RAND_116;
  reg [18:0] _T_117_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177651.4]
  reg [31:0] _RAND_117;
  reg [18:0] _T_118_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177656.4]
  reg [31:0] _RAND_118;
  reg [18:0] _T_119_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177661.4]
  reg [31:0] _RAND_119;
  reg [18:0] _T_120_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177666.4]
  reg [31:0] _RAND_120;
  reg [18:0] _T_121_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177671.4]
  reg [31:0] _RAND_121;
  reg [7:0] _T_122_0; // @[Mesh.scala 48:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@177676.4]
  reg [31:0] _RAND_122;
  reg  _T_123_0; // @[Mesh.scala 48:52:example.TestHarness.GemminiSocTest1RocketConfig.fir@177678.4]
  reg [31:0] _RAND_123;
  reg [7:0] _T_124_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177680.4]
  reg [31:0] _RAND_124;
  reg [18:0] _T_125_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177685.4]
  reg [31:0] _RAND_125;
  reg [18:0] _T_126_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177690.4]
  reg [31:0] _RAND_126;
  reg [18:0] _T_127_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177695.4]
  reg [31:0] _RAND_127;
  reg [18:0] _T_128_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177700.4]
  reg [31:0] _RAND_128;
  reg [18:0] _T_129_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177705.4]
  reg [31:0] _RAND_129;
  reg [18:0] _T_130_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177710.4]
  reg [31:0] _RAND_130;
  reg [18:0] _T_131_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177715.4]
  reg [31:0] _RAND_131;
  reg [7:0] _T_132_0; // @[Mesh.scala 48:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@177720.4]
  reg [31:0] _RAND_132;
  reg  _T_133_0; // @[Mesh.scala 48:52:example.TestHarness.GemminiSocTest1RocketConfig.fir@177722.4]
  reg [31:0] _RAND_133;
  reg [7:0] _T_134_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177724.4]
  reg [31:0] _RAND_134;
  reg [18:0] _T_135_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177729.4]
  reg [31:0] _RAND_135;
  reg [18:0] _T_136_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177734.4]
  reg [31:0] _RAND_136;
  reg [18:0] _T_137_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177739.4]
  reg [31:0] _RAND_137;
  reg [18:0] _T_138_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177744.4]
  reg [31:0] _RAND_138;
  reg [18:0] _T_139_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177749.4]
  reg [31:0] _RAND_139;
  reg [18:0] _T_140_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177754.4]
  reg [31:0] _RAND_140;
  reg [18:0] _T_141_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177759.4]
  reg [31:0] _RAND_141;
  reg [7:0] _T_142_0; // @[Mesh.scala 48:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@177764.4]
  reg [31:0] _RAND_142;
  reg  _T_143_0; // @[Mesh.scala 48:52:example.TestHarness.GemminiSocTest1RocketConfig.fir@177766.4]
  reg [31:0] _RAND_143;
  reg [7:0] _T_144_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177768.4]
  reg [31:0] _RAND_144;
  reg [18:0] _T_145_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177773.4]
  reg [31:0] _RAND_145;
  reg [18:0] _T_146_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177778.4]
  reg [31:0] _RAND_146;
  reg [18:0] _T_147_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177783.4]
  reg [31:0] _RAND_147;
  reg [18:0] _T_148_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177788.4]
  reg [31:0] _RAND_148;
  reg [18:0] _T_149_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177793.4]
  reg [31:0] _RAND_149;
  reg [18:0] _T_150_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177798.4]
  reg [31:0] _RAND_150;
  reg [18:0] _T_151_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177803.4]
  reg [31:0] _RAND_151;
  reg [7:0] _T_152_0; // @[Mesh.scala 56:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@177808.4]
  reg [31:0] _RAND_152;
  reg  _T_153_0; // @[Mesh.scala 56:52:example.TestHarness.GemminiSocTest1RocketConfig.fir@177810.4]
  reg [31:0] _RAND_153;
  reg [7:0] _T_154_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177812.4]
  reg [31:0] _RAND_154;
  reg [18:0] _T_155_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177817.4]
  reg [31:0] _RAND_155;
  reg [18:0] _T_156_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177822.4]
  reg [31:0] _RAND_156;
  reg [18:0] _T_157_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177827.4]
  reg [31:0] _RAND_157;
  reg [18:0] _T_158_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177832.4]
  reg [31:0] _RAND_158;
  reg [18:0] _T_159_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177837.4]
  reg [31:0] _RAND_159;
  reg [18:0] _T_160_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177842.4]
  reg [31:0] _RAND_160;
  reg [18:0] _T_161_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177847.4]
  reg [31:0] _RAND_161;
  reg [7:0] _T_162_0; // @[Mesh.scala 56:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@177852.4]
  reg [31:0] _RAND_162;
  reg  _T_163_0; // @[Mesh.scala 56:52:example.TestHarness.GemminiSocTest1RocketConfig.fir@177854.4]
  reg [31:0] _RAND_163;
  reg [7:0] _T_164_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177856.4]
  reg [31:0] _RAND_164;
  reg [18:0] _T_165_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177861.4]
  reg [31:0] _RAND_165;
  reg [18:0] _T_166_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177866.4]
  reg [31:0] _RAND_166;
  reg [18:0] _T_167_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177871.4]
  reg [31:0] _RAND_167;
  reg [18:0] _T_168_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177876.4]
  reg [31:0] _RAND_168;
  reg [18:0] _T_169_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177881.4]
  reg [31:0] _RAND_169;
  reg [18:0] _T_170_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177886.4]
  reg [31:0] _RAND_170;
  reg [18:0] _T_171_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177891.4]
  reg [31:0] _RAND_171;
  reg [7:0] _T_172_0; // @[Mesh.scala 56:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@177896.4]
  reg [31:0] _RAND_172;
  reg  _T_173_0; // @[Mesh.scala 56:52:example.TestHarness.GemminiSocTest1RocketConfig.fir@177898.4]
  reg [31:0] _RAND_173;
  reg [7:0] _T_174_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177900.4]
  reg [31:0] _RAND_174;
  reg [18:0] _T_175_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177905.4]
  reg [31:0] _RAND_175;
  reg [18:0] _T_176_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177910.4]
  reg [31:0] _RAND_176;
  reg [18:0] _T_177_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177915.4]
  reg [31:0] _RAND_177;
  reg [18:0] _T_178_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177920.4]
  reg [31:0] _RAND_178;
  reg [18:0] _T_179_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177925.4]
  reg [31:0] _RAND_179;
  reg [18:0] _T_180_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177930.4]
  reg [31:0] _RAND_180;
  reg [18:0] _T_181_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177935.4]
  reg [31:0] _RAND_181;
  reg [7:0] _T_182_0; // @[Mesh.scala 56:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@177940.4]
  reg [31:0] _RAND_182;
  reg  _T_183_0; // @[Mesh.scala 56:52:example.TestHarness.GemminiSocTest1RocketConfig.fir@177942.4]
  reg [31:0] _RAND_183;
  reg [7:0] _T_184_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177944.4]
  reg [31:0] _RAND_184;
  reg [18:0] _T_185_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177949.4]
  reg [31:0] _RAND_185;
  reg [18:0] _T_186_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177954.4]
  reg [31:0] _RAND_186;
  reg [18:0] _T_187_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177959.4]
  reg [31:0] _RAND_187;
  reg [18:0] _T_188_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177964.4]
  reg [31:0] _RAND_188;
  reg [18:0] _T_189_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177969.4]
  reg [31:0] _RAND_189;
  reg [18:0] _T_190_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177974.4]
  reg [31:0] _RAND_190;
  reg [18:0] _T_191_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177979.4]
  reg [31:0] _RAND_191;
  reg [7:0] _T_192_0; // @[Mesh.scala 56:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@177984.4]
  reg [31:0] _RAND_192;
  reg  _T_193_0; // @[Mesh.scala 56:52:example.TestHarness.GemminiSocTest1RocketConfig.fir@177986.4]
  reg [31:0] _RAND_193;
  reg [7:0] _T_194_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177988.4]
  reg [31:0] _RAND_194;
  reg [18:0] _T_195_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177993.4]
  reg [31:0] _RAND_195;
  reg [18:0] _T_196_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@177998.4]
  reg [31:0] _RAND_196;
  reg [18:0] _T_197_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178003.4]
  reg [31:0] _RAND_197;
  reg [18:0] _T_198_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178008.4]
  reg [31:0] _RAND_198;
  reg [18:0] _T_199_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178013.4]
  reg [31:0] _RAND_199;
  reg [18:0] _T_200_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178018.4]
  reg [31:0] _RAND_200;
  reg [18:0] _T_201_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178023.4]
  reg [31:0] _RAND_201;
  reg [7:0] _T_202_0; // @[Mesh.scala 56:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178028.4]
  reg [31:0] _RAND_202;
  reg  _T_203_0; // @[Mesh.scala 56:52:example.TestHarness.GemminiSocTest1RocketConfig.fir@178030.4]
  reg [31:0] _RAND_203;
  reg [7:0] _T_204_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178032.4]
  reg [31:0] _RAND_204;
  reg [18:0] _T_205_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178037.4]
  reg [31:0] _RAND_205;
  reg [18:0] _T_206_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178042.4]
  reg [31:0] _RAND_206;
  reg [18:0] _T_207_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178047.4]
  reg [31:0] _RAND_207;
  reg [18:0] _T_208_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178052.4]
  reg [31:0] _RAND_208;
  reg [18:0] _T_209_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178057.4]
  reg [31:0] _RAND_209;
  reg [18:0] _T_210_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178062.4]
  reg [31:0] _RAND_210;
  reg [18:0] _T_211_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178067.4]
  reg [31:0] _RAND_211;
  reg [7:0] _T_212_0; // @[Mesh.scala 56:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178072.4]
  reg [31:0] _RAND_212;
  reg  _T_213_0; // @[Mesh.scala 56:52:example.TestHarness.GemminiSocTest1RocketConfig.fir@178074.4]
  reg [31:0] _RAND_213;
  reg [7:0] _T_214_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178076.4]
  reg [31:0] _RAND_214;
  reg [18:0] _T_215_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178081.4]
  reg [31:0] _RAND_215;
  reg [18:0] _T_216_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178086.4]
  reg [31:0] _RAND_216;
  reg [18:0] _T_217_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178091.4]
  reg [31:0] _RAND_217;
  reg [18:0] _T_218_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178096.4]
  reg [31:0] _RAND_218;
  reg [18:0] _T_219_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178101.4]
  reg [31:0] _RAND_219;
  reg [18:0] _T_220_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178106.4]
  reg [31:0] _RAND_220;
  reg [18:0] _T_221_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178111.4]
  reg [31:0] _RAND_221;
  reg [7:0] _T_222_0; // @[Mesh.scala 56:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178116.4]
  reg [31:0] _RAND_222;
  reg  _T_223_0; // @[Mesh.scala 56:52:example.TestHarness.GemminiSocTest1RocketConfig.fir@178118.4]
  reg [31:0] _RAND_223;
  reg [7:0] _T_224_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178120.4]
  reg [31:0] _RAND_224;
  reg [18:0] _T_225_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178125.4]
  reg [31:0] _RAND_225;
  reg [18:0] _T_226_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178130.4]
  reg [31:0] _RAND_226;
  reg [18:0] _T_227_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178135.4]
  reg [31:0] _RAND_227;
  reg [18:0] _T_228_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178140.4]
  reg [31:0] _RAND_228;
  reg [18:0] _T_229_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178145.4]
  reg [31:0] _RAND_229;
  reg [18:0] _T_230_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178150.4]
  reg [31:0] _RAND_230;
  reg [18:0] _T_231_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178155.4]
  reg [31:0] _RAND_231;
  reg  _T_232_0_propagate; // @[Mesh.scala 64:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178160.4]
  reg [31:0] _RAND_232;
  reg [4:0] _T_232_0_shift; // @[Mesh.scala 64:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178160.4]
  reg [31:0] _RAND_233;
  reg  _T_233_0; // @[Mesh.scala 64:58:example.TestHarness.GemminiSocTest1RocketConfig.fir@178164.4]
  reg [31:0] _RAND_234;
  reg [4:0] _T_234; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178166.4]
  reg [31:0] _RAND_235;
  reg  _T_236; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178176.4]
  reg [31:0] _RAND_236;
  reg [4:0] _T_237; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178181.4]
  reg [31:0] _RAND_237;
  reg  _T_239; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178191.4]
  reg [31:0] _RAND_238;
  reg [4:0] _T_240; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178196.4]
  reg [31:0] _RAND_239;
  reg  _T_242; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178206.4]
  reg [31:0] _RAND_240;
  reg [4:0] _T_243; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178211.4]
  reg [31:0] _RAND_241;
  reg  _T_245; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178221.4]
  reg [31:0] _RAND_242;
  reg [4:0] _T_246; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178226.4]
  reg [31:0] _RAND_243;
  reg  _T_248; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178236.4]
  reg [31:0] _RAND_244;
  reg [4:0] _T_249; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178241.4]
  reg [31:0] _RAND_245;
  reg  _T_251; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178251.4]
  reg [31:0] _RAND_246;
  reg [4:0] _T_252; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178256.4]
  reg [31:0] _RAND_247;
  reg  _T_254; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178266.4]
  reg [31:0] _RAND_248;
  reg [4:0] _T_255; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178271.4]
  reg [31:0] _RAND_249;
  reg  _T_257; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178281.4]
  reg [31:0] _RAND_250;
  reg  _T_258_0_propagate; // @[Mesh.scala 64:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178286.4]
  reg [31:0] _RAND_251;
  reg [4:0] _T_258_0_shift; // @[Mesh.scala 64:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178286.4]
  reg [31:0] _RAND_252;
  reg  _T_259_0; // @[Mesh.scala 64:58:example.TestHarness.GemminiSocTest1RocketConfig.fir@178290.4]
  reg [31:0] _RAND_253;
  reg [4:0] _T_260; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178292.4]
  reg [31:0] _RAND_254;
  reg  _T_262; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178302.4]
  reg [31:0] _RAND_255;
  reg [4:0] _T_263; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178307.4]
  reg [31:0] _RAND_256;
  reg  _T_265; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178317.4]
  reg [31:0] _RAND_257;
  reg [4:0] _T_266; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178322.4]
  reg [31:0] _RAND_258;
  reg  _T_268; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178332.4]
  reg [31:0] _RAND_259;
  reg [4:0] _T_269; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178337.4]
  reg [31:0] _RAND_260;
  reg  _T_271; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178347.4]
  reg [31:0] _RAND_261;
  reg [4:0] _T_272; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178352.4]
  reg [31:0] _RAND_262;
  reg  _T_274; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178362.4]
  reg [31:0] _RAND_263;
  reg [4:0] _T_275; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178367.4]
  reg [31:0] _RAND_264;
  reg  _T_277; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178377.4]
  reg [31:0] _RAND_265;
  reg [4:0] _T_278; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178382.4]
  reg [31:0] _RAND_266;
  reg  _T_280; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178392.4]
  reg [31:0] _RAND_267;
  reg [4:0] _T_281; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178397.4]
  reg [31:0] _RAND_268;
  reg  _T_283; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178407.4]
  reg [31:0] _RAND_269;
  reg  _T_284_0_propagate; // @[Mesh.scala 64:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178412.4]
  reg [31:0] _RAND_270;
  reg [4:0] _T_284_0_shift; // @[Mesh.scala 64:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178412.4]
  reg [31:0] _RAND_271;
  reg  _T_285_0; // @[Mesh.scala 64:58:example.TestHarness.GemminiSocTest1RocketConfig.fir@178416.4]
  reg [31:0] _RAND_272;
  reg [4:0] _T_286; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178418.4]
  reg [31:0] _RAND_273;
  reg  _T_288; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178428.4]
  reg [31:0] _RAND_274;
  reg [4:0] _T_289; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178433.4]
  reg [31:0] _RAND_275;
  reg  _T_291; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178443.4]
  reg [31:0] _RAND_276;
  reg [4:0] _T_292; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178448.4]
  reg [31:0] _RAND_277;
  reg  _T_294; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178458.4]
  reg [31:0] _RAND_278;
  reg [4:0] _T_295; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178463.4]
  reg [31:0] _RAND_279;
  reg  _T_297; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178473.4]
  reg [31:0] _RAND_280;
  reg [4:0] _T_298; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178478.4]
  reg [31:0] _RAND_281;
  reg  _T_300; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178488.4]
  reg [31:0] _RAND_282;
  reg [4:0] _T_301; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178493.4]
  reg [31:0] _RAND_283;
  reg  _T_303; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178503.4]
  reg [31:0] _RAND_284;
  reg [4:0] _T_304; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178508.4]
  reg [31:0] _RAND_285;
  reg  _T_306; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178518.4]
  reg [31:0] _RAND_286;
  reg [4:0] _T_307; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178523.4]
  reg [31:0] _RAND_287;
  reg  _T_309; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178533.4]
  reg [31:0] _RAND_288;
  reg  _T_310_0_propagate; // @[Mesh.scala 64:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178538.4]
  reg [31:0] _RAND_289;
  reg [4:0] _T_310_0_shift; // @[Mesh.scala 64:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178538.4]
  reg [31:0] _RAND_290;
  reg  _T_311_0; // @[Mesh.scala 64:58:example.TestHarness.GemminiSocTest1RocketConfig.fir@178542.4]
  reg [31:0] _RAND_291;
  reg [4:0] _T_312; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178544.4]
  reg [31:0] _RAND_292;
  reg  _T_314; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178554.4]
  reg [31:0] _RAND_293;
  reg [4:0] _T_315; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178559.4]
  reg [31:0] _RAND_294;
  reg  _T_317; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178569.4]
  reg [31:0] _RAND_295;
  reg [4:0] _T_318; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178574.4]
  reg [31:0] _RAND_296;
  reg  _T_320; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178584.4]
  reg [31:0] _RAND_297;
  reg [4:0] _T_321; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178589.4]
  reg [31:0] _RAND_298;
  reg  _T_323; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178599.4]
  reg [31:0] _RAND_299;
  reg [4:0] _T_324; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178604.4]
  reg [31:0] _RAND_300;
  reg  _T_326; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178614.4]
  reg [31:0] _RAND_301;
  reg [4:0] _T_327; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178619.4]
  reg [31:0] _RAND_302;
  reg  _T_329; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178629.4]
  reg [31:0] _RAND_303;
  reg [4:0] _T_330; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178634.4]
  reg [31:0] _RAND_304;
  reg  _T_332; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178644.4]
  reg [31:0] _RAND_305;
  reg [4:0] _T_333; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178649.4]
  reg [31:0] _RAND_306;
  reg  _T_335; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178659.4]
  reg [31:0] _RAND_307;
  reg  _T_336_0_propagate; // @[Mesh.scala 64:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178664.4]
  reg [31:0] _RAND_308;
  reg [4:0] _T_336_0_shift; // @[Mesh.scala 64:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178664.4]
  reg [31:0] _RAND_309;
  reg  _T_337_0; // @[Mesh.scala 64:58:example.TestHarness.GemminiSocTest1RocketConfig.fir@178668.4]
  reg [31:0] _RAND_310;
  reg [4:0] _T_338; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178670.4]
  reg [31:0] _RAND_311;
  reg  _T_340; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178680.4]
  reg [31:0] _RAND_312;
  reg [4:0] _T_341; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178685.4]
  reg [31:0] _RAND_313;
  reg  _T_343; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178695.4]
  reg [31:0] _RAND_314;
  reg [4:0] _T_344; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178700.4]
  reg [31:0] _RAND_315;
  reg  _T_346; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178710.4]
  reg [31:0] _RAND_316;
  reg [4:0] _T_347; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178715.4]
  reg [31:0] _RAND_317;
  reg  _T_349; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178725.4]
  reg [31:0] _RAND_318;
  reg [4:0] _T_350; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178730.4]
  reg [31:0] _RAND_319;
  reg  _T_352; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178740.4]
  reg [31:0] _RAND_320;
  reg [4:0] _T_353; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178745.4]
  reg [31:0] _RAND_321;
  reg  _T_355; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178755.4]
  reg [31:0] _RAND_322;
  reg [4:0] _T_356; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178760.4]
  reg [31:0] _RAND_323;
  reg  _T_358; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178770.4]
  reg [31:0] _RAND_324;
  reg [4:0] _T_359; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178775.4]
  reg [31:0] _RAND_325;
  reg  _T_361; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178785.4]
  reg [31:0] _RAND_326;
  reg  _T_362_0_propagate; // @[Mesh.scala 64:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178790.4]
  reg [31:0] _RAND_327;
  reg [4:0] _T_362_0_shift; // @[Mesh.scala 64:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178790.4]
  reg [31:0] _RAND_328;
  reg  _T_363_0; // @[Mesh.scala 64:58:example.TestHarness.GemminiSocTest1RocketConfig.fir@178794.4]
  reg [31:0] _RAND_329;
  reg [4:0] _T_364; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178796.4]
  reg [31:0] _RAND_330;
  reg  _T_366; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178806.4]
  reg [31:0] _RAND_331;
  reg [4:0] _T_367; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178811.4]
  reg [31:0] _RAND_332;
  reg  _T_369; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178821.4]
  reg [31:0] _RAND_333;
  reg [4:0] _T_370; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178826.4]
  reg [31:0] _RAND_334;
  reg  _T_372; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178836.4]
  reg [31:0] _RAND_335;
  reg [4:0] _T_373; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178841.4]
  reg [31:0] _RAND_336;
  reg  _T_375; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178851.4]
  reg [31:0] _RAND_337;
  reg [4:0] _T_376; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178856.4]
  reg [31:0] _RAND_338;
  reg  _T_378; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178866.4]
  reg [31:0] _RAND_339;
  reg [4:0] _T_379; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178871.4]
  reg [31:0] _RAND_340;
  reg  _T_381; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178881.4]
  reg [31:0] _RAND_341;
  reg [4:0] _T_382; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178886.4]
  reg [31:0] _RAND_342;
  reg  _T_384; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178896.4]
  reg [31:0] _RAND_343;
  reg [4:0] _T_385; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178901.4]
  reg [31:0] _RAND_344;
  reg  _T_387; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178911.4]
  reg [31:0] _RAND_345;
  reg  _T_388_0_propagate; // @[Mesh.scala 64:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178916.4]
  reg [31:0] _RAND_346;
  reg [4:0] _T_388_0_shift; // @[Mesh.scala 64:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178916.4]
  reg [31:0] _RAND_347;
  reg  _T_389_0; // @[Mesh.scala 64:58:example.TestHarness.GemminiSocTest1RocketConfig.fir@178920.4]
  reg [31:0] _RAND_348;
  reg [4:0] _T_390; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178922.4]
  reg [31:0] _RAND_349;
  reg  _T_392; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178932.4]
  reg [31:0] _RAND_350;
  reg [4:0] _T_393; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178937.4]
  reg [31:0] _RAND_351;
  reg  _T_395; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178947.4]
  reg [31:0] _RAND_352;
  reg [4:0] _T_396; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178952.4]
  reg [31:0] _RAND_353;
  reg  _T_398; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178962.4]
  reg [31:0] _RAND_354;
  reg [4:0] _T_399; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178967.4]
  reg [31:0] _RAND_355;
  reg  _T_401; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178977.4]
  reg [31:0] _RAND_356;
  reg [4:0] _T_402; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178982.4]
  reg [31:0] _RAND_357;
  reg  _T_404; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178992.4]
  reg [31:0] _RAND_358;
  reg [4:0] _T_405; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@178997.4]
  reg [31:0] _RAND_359;
  reg  _T_407; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@179007.4]
  reg [31:0] _RAND_360;
  reg [4:0] _T_408; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@179012.4]
  reg [31:0] _RAND_361;
  reg  _T_410; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@179022.4]
  reg [31:0] _RAND_362;
  reg [4:0] _T_411; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@179027.4]
  reg [31:0] _RAND_363;
  reg  _T_413; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@179037.4]
  reg [31:0] _RAND_364;
  reg  _T_414_0_propagate; // @[Mesh.scala 64:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@179042.4]
  reg [31:0] _RAND_365;
  reg [4:0] _T_414_0_shift; // @[Mesh.scala 64:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@179042.4]
  reg [31:0] _RAND_366;
  reg  _T_415_0; // @[Mesh.scala 64:58:example.TestHarness.GemminiSocTest1RocketConfig.fir@179046.4]
  reg [31:0] _RAND_367;
  reg [4:0] _T_416; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@179048.4]
  reg [31:0] _RAND_368;
  reg  _T_418; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@179058.4]
  reg [31:0] _RAND_369;
  reg [4:0] _T_419; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@179063.4]
  reg [31:0] _RAND_370;
  reg  _T_421; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@179073.4]
  reg [31:0] _RAND_371;
  reg [4:0] _T_422; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@179078.4]
  reg [31:0] _RAND_372;
  reg  _T_424; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@179088.4]
  reg [31:0] _RAND_373;
  reg [4:0] _T_425; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@179093.4]
  reg [31:0] _RAND_374;
  reg  _T_427; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@179103.4]
  reg [31:0] _RAND_375;
  reg [4:0] _T_428; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@179108.4]
  reg [31:0] _RAND_376;
  reg  _T_430; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@179118.4]
  reg [31:0] _RAND_377;
  reg [4:0] _T_431; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@179123.4]
  reg [31:0] _RAND_378;
  reg  _T_433; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@179133.4]
  reg [31:0] _RAND_379;
  reg [4:0] _T_434; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@179138.4]
  reg [31:0] _RAND_380;
  reg  _T_436; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@179148.4]
  reg [31:0] _RAND_381;
  reg [4:0] _T_437; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@179153.4]
  reg [31:0] _RAND_382;
  reg  _T_439; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig.fir@179163.4]
  reg [31:0] _RAND_383;
  reg  _T_440_0; // @[Mesh.scala 76:30:example.TestHarness.GemminiSocTest1RocketConfig.fir@179168.4]
  reg [31:0] _RAND_384;
  reg  _T_441_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179170.4]
  reg [31:0] _RAND_385;
  reg  _T_442_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179173.4]
  reg [31:0] _RAND_386;
  reg  _T_443_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179176.4]
  reg [31:0] _RAND_387;
  reg  _T_444_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179179.4]
  reg [31:0] _RAND_388;
  reg  _T_445_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179182.4]
  reg [31:0] _RAND_389;
  reg  _T_446_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179185.4]
  reg [31:0] _RAND_390;
  reg  _T_447_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179188.4]
  reg [31:0] _RAND_391;
  reg  _T_448_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179191.4]
  reg [31:0] _RAND_392;
  reg  _T_449_0; // @[Mesh.scala 76:30:example.TestHarness.GemminiSocTest1RocketConfig.fir@179194.4]
  reg [31:0] _RAND_393;
  reg  _T_450_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179196.4]
  reg [31:0] _RAND_394;
  reg  _T_451_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179199.4]
  reg [31:0] _RAND_395;
  reg  _T_452_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179202.4]
  reg [31:0] _RAND_396;
  reg  _T_453_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179205.4]
  reg [31:0] _RAND_397;
  reg  _T_454_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179208.4]
  reg [31:0] _RAND_398;
  reg  _T_455_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179211.4]
  reg [31:0] _RAND_399;
  reg  _T_456_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179214.4]
  reg [31:0] _RAND_400;
  reg  _T_457_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179217.4]
  reg [31:0] _RAND_401;
  reg  _T_458_0; // @[Mesh.scala 76:30:example.TestHarness.GemminiSocTest1RocketConfig.fir@179220.4]
  reg [31:0] _RAND_402;
  reg  _T_459_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179222.4]
  reg [31:0] _RAND_403;
  reg  _T_460_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179225.4]
  reg [31:0] _RAND_404;
  reg  _T_461_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179228.4]
  reg [31:0] _RAND_405;
  reg  _T_462_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179231.4]
  reg [31:0] _RAND_406;
  reg  _T_463_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179234.4]
  reg [31:0] _RAND_407;
  reg  _T_464_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179237.4]
  reg [31:0] _RAND_408;
  reg  _T_465_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179240.4]
  reg [31:0] _RAND_409;
  reg  _T_466_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179243.4]
  reg [31:0] _RAND_410;
  reg  _T_467_0; // @[Mesh.scala 76:30:example.TestHarness.GemminiSocTest1RocketConfig.fir@179246.4]
  reg [31:0] _RAND_411;
  reg  _T_468_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179248.4]
  reg [31:0] _RAND_412;
  reg  _T_469_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179251.4]
  reg [31:0] _RAND_413;
  reg  _T_470_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179254.4]
  reg [31:0] _RAND_414;
  reg  _T_471_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179257.4]
  reg [31:0] _RAND_415;
  reg  _T_472_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179260.4]
  reg [31:0] _RAND_416;
  reg  _T_473_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179263.4]
  reg [31:0] _RAND_417;
  reg  _T_474_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179266.4]
  reg [31:0] _RAND_418;
  reg  _T_475_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179269.4]
  reg [31:0] _RAND_419;
  reg  _T_476_0; // @[Mesh.scala 76:30:example.TestHarness.GemminiSocTest1RocketConfig.fir@179272.4]
  reg [31:0] _RAND_420;
  reg  _T_477_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179274.4]
  reg [31:0] _RAND_421;
  reg  _T_478_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179277.4]
  reg [31:0] _RAND_422;
  reg  _T_479_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179280.4]
  reg [31:0] _RAND_423;
  reg  _T_480_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179283.4]
  reg [31:0] _RAND_424;
  reg  _T_481_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179286.4]
  reg [31:0] _RAND_425;
  reg  _T_482_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179289.4]
  reg [31:0] _RAND_426;
  reg  _T_483_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179292.4]
  reg [31:0] _RAND_427;
  reg  _T_484_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179295.4]
  reg [31:0] _RAND_428;
  reg  _T_485_0; // @[Mesh.scala 76:30:example.TestHarness.GemminiSocTest1RocketConfig.fir@179298.4]
  reg [31:0] _RAND_429;
  reg  _T_486_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179300.4]
  reg [31:0] _RAND_430;
  reg  _T_487_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179303.4]
  reg [31:0] _RAND_431;
  reg  _T_488_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179306.4]
  reg [31:0] _RAND_432;
  reg  _T_489_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179309.4]
  reg [31:0] _RAND_433;
  reg  _T_490_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179312.4]
  reg [31:0] _RAND_434;
  reg  _T_491_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179315.4]
  reg [31:0] _RAND_435;
  reg  _T_492_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179318.4]
  reg [31:0] _RAND_436;
  reg  _T_493_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179321.4]
  reg [31:0] _RAND_437;
  reg  _T_494_0; // @[Mesh.scala 76:30:example.TestHarness.GemminiSocTest1RocketConfig.fir@179324.4]
  reg [31:0] _RAND_438;
  reg  _T_495_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179326.4]
  reg [31:0] _RAND_439;
  reg  _T_496_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179329.4]
  reg [31:0] _RAND_440;
  reg  _T_497_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179332.4]
  reg [31:0] _RAND_441;
  reg  _T_498_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179335.4]
  reg [31:0] _RAND_442;
  reg  _T_499_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179338.4]
  reg [31:0] _RAND_443;
  reg  _T_500_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179341.4]
  reg [31:0] _RAND_444;
  reg  _T_501_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179344.4]
  reg [31:0] _RAND_445;
  reg  _T_502_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179347.4]
  reg [31:0] _RAND_446;
  reg  _T_503_0; // @[Mesh.scala 76:30:example.TestHarness.GemminiSocTest1RocketConfig.fir@179350.4]
  reg [31:0] _RAND_447;
  reg  _T_504_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179352.4]
  reg [31:0] _RAND_448;
  reg  _T_505_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179355.4]
  reg [31:0] _RAND_449;
  reg  _T_506_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179358.4]
  reg [31:0] _RAND_450;
  reg  _T_507_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179361.4]
  reg [31:0] _RAND_451;
  reg  _T_508_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179364.4]
  reg [31:0] _RAND_452;
  reg  _T_509_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179367.4]
  reg [31:0] _RAND_453;
  reg  _T_510_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179370.4]
  reg [31:0] _RAND_454;
  reg  _T_511_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig.fir@179373.4]
  reg [31:0] _RAND_455;
  Tile mesh_0_0 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177056.4]
    .clock(mesh_0_0_clock),
    .io_in_a_0(mesh_0_0_io_in_a_0),
    .io_in_b_0(mesh_0_0_io_in_b_0),
    .io_in_d_0(mesh_0_0_io_in_d_0),
    .io_in_control_0_propagate(mesh_0_0_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_0_0_io_in_control_0_shift),
    .io_out_a_0(mesh_0_0_io_out_a_0),
    .io_out_c_0(mesh_0_0_io_out_c_0),
    .io_out_b_0(mesh_0_0_io_out_b_0),
    .io_out_control_0_propagate(mesh_0_0_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_0_0_io_out_control_0_shift),
    .io_in_valid_0(mesh_0_0_io_in_valid_0),
    .io_out_valid_0(mesh_0_0_io_out_valid_0)
  );
  Tile mesh_0_1 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177059.4]
    .clock(mesh_0_1_clock),
    .io_in_a_0(mesh_0_1_io_in_a_0),
    .io_in_b_0(mesh_0_1_io_in_b_0),
    .io_in_d_0(mesh_0_1_io_in_d_0),
    .io_in_control_0_propagate(mesh_0_1_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_0_1_io_in_control_0_shift),
    .io_out_a_0(mesh_0_1_io_out_a_0),
    .io_out_c_0(mesh_0_1_io_out_c_0),
    .io_out_b_0(mesh_0_1_io_out_b_0),
    .io_out_control_0_propagate(mesh_0_1_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_0_1_io_out_control_0_shift),
    .io_in_valid_0(mesh_0_1_io_in_valid_0),
    .io_out_valid_0(mesh_0_1_io_out_valid_0)
  );
  Tile mesh_0_2 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177062.4]
    .clock(mesh_0_2_clock),
    .io_in_a_0(mesh_0_2_io_in_a_0),
    .io_in_b_0(mesh_0_2_io_in_b_0),
    .io_in_d_0(mesh_0_2_io_in_d_0),
    .io_in_control_0_propagate(mesh_0_2_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_0_2_io_in_control_0_shift),
    .io_out_a_0(mesh_0_2_io_out_a_0),
    .io_out_c_0(mesh_0_2_io_out_c_0),
    .io_out_b_0(mesh_0_2_io_out_b_0),
    .io_out_control_0_propagate(mesh_0_2_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_0_2_io_out_control_0_shift),
    .io_in_valid_0(mesh_0_2_io_in_valid_0),
    .io_out_valid_0(mesh_0_2_io_out_valid_0)
  );
  Tile mesh_0_3 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177065.4]
    .clock(mesh_0_3_clock),
    .io_in_a_0(mesh_0_3_io_in_a_0),
    .io_in_b_0(mesh_0_3_io_in_b_0),
    .io_in_d_0(mesh_0_3_io_in_d_0),
    .io_in_control_0_propagate(mesh_0_3_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_0_3_io_in_control_0_shift),
    .io_out_a_0(mesh_0_3_io_out_a_0),
    .io_out_c_0(mesh_0_3_io_out_c_0),
    .io_out_b_0(mesh_0_3_io_out_b_0),
    .io_out_control_0_propagate(mesh_0_3_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_0_3_io_out_control_0_shift),
    .io_in_valid_0(mesh_0_3_io_in_valid_0),
    .io_out_valid_0(mesh_0_3_io_out_valid_0)
  );
  Tile mesh_0_4 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177068.4]
    .clock(mesh_0_4_clock),
    .io_in_a_0(mesh_0_4_io_in_a_0),
    .io_in_b_0(mesh_0_4_io_in_b_0),
    .io_in_d_0(mesh_0_4_io_in_d_0),
    .io_in_control_0_propagate(mesh_0_4_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_0_4_io_in_control_0_shift),
    .io_out_a_0(mesh_0_4_io_out_a_0),
    .io_out_c_0(mesh_0_4_io_out_c_0),
    .io_out_b_0(mesh_0_4_io_out_b_0),
    .io_out_control_0_propagate(mesh_0_4_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_0_4_io_out_control_0_shift),
    .io_in_valid_0(mesh_0_4_io_in_valid_0),
    .io_out_valid_0(mesh_0_4_io_out_valid_0)
  );
  Tile mesh_0_5 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177071.4]
    .clock(mesh_0_5_clock),
    .io_in_a_0(mesh_0_5_io_in_a_0),
    .io_in_b_0(mesh_0_5_io_in_b_0),
    .io_in_d_0(mesh_0_5_io_in_d_0),
    .io_in_control_0_propagate(mesh_0_5_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_0_5_io_in_control_0_shift),
    .io_out_a_0(mesh_0_5_io_out_a_0),
    .io_out_c_0(mesh_0_5_io_out_c_0),
    .io_out_b_0(mesh_0_5_io_out_b_0),
    .io_out_control_0_propagate(mesh_0_5_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_0_5_io_out_control_0_shift),
    .io_in_valid_0(mesh_0_5_io_in_valid_0),
    .io_out_valid_0(mesh_0_5_io_out_valid_0)
  );
  Tile mesh_0_6 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177074.4]
    .clock(mesh_0_6_clock),
    .io_in_a_0(mesh_0_6_io_in_a_0),
    .io_in_b_0(mesh_0_6_io_in_b_0),
    .io_in_d_0(mesh_0_6_io_in_d_0),
    .io_in_control_0_propagate(mesh_0_6_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_0_6_io_in_control_0_shift),
    .io_out_a_0(mesh_0_6_io_out_a_0),
    .io_out_c_0(mesh_0_6_io_out_c_0),
    .io_out_b_0(mesh_0_6_io_out_b_0),
    .io_out_control_0_propagate(mesh_0_6_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_0_6_io_out_control_0_shift),
    .io_in_valid_0(mesh_0_6_io_in_valid_0),
    .io_out_valid_0(mesh_0_6_io_out_valid_0)
  );
  Tile mesh_0_7 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177077.4]
    .clock(mesh_0_7_clock),
    .io_in_a_0(mesh_0_7_io_in_a_0),
    .io_in_b_0(mesh_0_7_io_in_b_0),
    .io_in_d_0(mesh_0_7_io_in_d_0),
    .io_in_control_0_propagate(mesh_0_7_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_0_7_io_in_control_0_shift),
    .io_out_a_0(mesh_0_7_io_out_a_0),
    .io_out_c_0(mesh_0_7_io_out_c_0),
    .io_out_b_0(mesh_0_7_io_out_b_0),
    .io_out_control_0_propagate(mesh_0_7_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_0_7_io_out_control_0_shift),
    .io_in_valid_0(mesh_0_7_io_in_valid_0),
    .io_out_valid_0(mesh_0_7_io_out_valid_0)
  );
  Tile mesh_1_0 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177080.4]
    .clock(mesh_1_0_clock),
    .io_in_a_0(mesh_1_0_io_in_a_0),
    .io_in_b_0(mesh_1_0_io_in_b_0),
    .io_in_d_0(mesh_1_0_io_in_d_0),
    .io_in_control_0_propagate(mesh_1_0_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_1_0_io_in_control_0_shift),
    .io_out_a_0(mesh_1_0_io_out_a_0),
    .io_out_c_0(mesh_1_0_io_out_c_0),
    .io_out_b_0(mesh_1_0_io_out_b_0),
    .io_out_control_0_propagate(mesh_1_0_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_1_0_io_out_control_0_shift),
    .io_in_valid_0(mesh_1_0_io_in_valid_0),
    .io_out_valid_0(mesh_1_0_io_out_valid_0)
  );
  Tile mesh_1_1 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177083.4]
    .clock(mesh_1_1_clock),
    .io_in_a_0(mesh_1_1_io_in_a_0),
    .io_in_b_0(mesh_1_1_io_in_b_0),
    .io_in_d_0(mesh_1_1_io_in_d_0),
    .io_in_control_0_propagate(mesh_1_1_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_1_1_io_in_control_0_shift),
    .io_out_a_0(mesh_1_1_io_out_a_0),
    .io_out_c_0(mesh_1_1_io_out_c_0),
    .io_out_b_0(mesh_1_1_io_out_b_0),
    .io_out_control_0_propagate(mesh_1_1_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_1_1_io_out_control_0_shift),
    .io_in_valid_0(mesh_1_1_io_in_valid_0),
    .io_out_valid_0(mesh_1_1_io_out_valid_0)
  );
  Tile mesh_1_2 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177086.4]
    .clock(mesh_1_2_clock),
    .io_in_a_0(mesh_1_2_io_in_a_0),
    .io_in_b_0(mesh_1_2_io_in_b_0),
    .io_in_d_0(mesh_1_2_io_in_d_0),
    .io_in_control_0_propagate(mesh_1_2_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_1_2_io_in_control_0_shift),
    .io_out_a_0(mesh_1_2_io_out_a_0),
    .io_out_c_0(mesh_1_2_io_out_c_0),
    .io_out_b_0(mesh_1_2_io_out_b_0),
    .io_out_control_0_propagate(mesh_1_2_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_1_2_io_out_control_0_shift),
    .io_in_valid_0(mesh_1_2_io_in_valid_0),
    .io_out_valid_0(mesh_1_2_io_out_valid_0)
  );
  Tile mesh_1_3 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177089.4]
    .clock(mesh_1_3_clock),
    .io_in_a_0(mesh_1_3_io_in_a_0),
    .io_in_b_0(mesh_1_3_io_in_b_0),
    .io_in_d_0(mesh_1_3_io_in_d_0),
    .io_in_control_0_propagate(mesh_1_3_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_1_3_io_in_control_0_shift),
    .io_out_a_0(mesh_1_3_io_out_a_0),
    .io_out_c_0(mesh_1_3_io_out_c_0),
    .io_out_b_0(mesh_1_3_io_out_b_0),
    .io_out_control_0_propagate(mesh_1_3_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_1_3_io_out_control_0_shift),
    .io_in_valid_0(mesh_1_3_io_in_valid_0),
    .io_out_valid_0(mesh_1_3_io_out_valid_0)
  );
  Tile mesh_1_4 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177092.4]
    .clock(mesh_1_4_clock),
    .io_in_a_0(mesh_1_4_io_in_a_0),
    .io_in_b_0(mesh_1_4_io_in_b_0),
    .io_in_d_0(mesh_1_4_io_in_d_0),
    .io_in_control_0_propagate(mesh_1_4_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_1_4_io_in_control_0_shift),
    .io_out_a_0(mesh_1_4_io_out_a_0),
    .io_out_c_0(mesh_1_4_io_out_c_0),
    .io_out_b_0(mesh_1_4_io_out_b_0),
    .io_out_control_0_propagate(mesh_1_4_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_1_4_io_out_control_0_shift),
    .io_in_valid_0(mesh_1_4_io_in_valid_0),
    .io_out_valid_0(mesh_1_4_io_out_valid_0)
  );
  Tile mesh_1_5 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177095.4]
    .clock(mesh_1_5_clock),
    .io_in_a_0(mesh_1_5_io_in_a_0),
    .io_in_b_0(mesh_1_5_io_in_b_0),
    .io_in_d_0(mesh_1_5_io_in_d_0),
    .io_in_control_0_propagate(mesh_1_5_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_1_5_io_in_control_0_shift),
    .io_out_a_0(mesh_1_5_io_out_a_0),
    .io_out_c_0(mesh_1_5_io_out_c_0),
    .io_out_b_0(mesh_1_5_io_out_b_0),
    .io_out_control_0_propagate(mesh_1_5_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_1_5_io_out_control_0_shift),
    .io_in_valid_0(mesh_1_5_io_in_valid_0),
    .io_out_valid_0(mesh_1_5_io_out_valid_0)
  );
  Tile mesh_1_6 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177098.4]
    .clock(mesh_1_6_clock),
    .io_in_a_0(mesh_1_6_io_in_a_0),
    .io_in_b_0(mesh_1_6_io_in_b_0),
    .io_in_d_0(mesh_1_6_io_in_d_0),
    .io_in_control_0_propagate(mesh_1_6_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_1_6_io_in_control_0_shift),
    .io_out_a_0(mesh_1_6_io_out_a_0),
    .io_out_c_0(mesh_1_6_io_out_c_0),
    .io_out_b_0(mesh_1_6_io_out_b_0),
    .io_out_control_0_propagate(mesh_1_6_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_1_6_io_out_control_0_shift),
    .io_in_valid_0(mesh_1_6_io_in_valid_0),
    .io_out_valid_0(mesh_1_6_io_out_valid_0)
  );
  Tile mesh_1_7 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177101.4]
    .clock(mesh_1_7_clock),
    .io_in_a_0(mesh_1_7_io_in_a_0),
    .io_in_b_0(mesh_1_7_io_in_b_0),
    .io_in_d_0(mesh_1_7_io_in_d_0),
    .io_in_control_0_propagate(mesh_1_7_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_1_7_io_in_control_0_shift),
    .io_out_a_0(mesh_1_7_io_out_a_0),
    .io_out_c_0(mesh_1_7_io_out_c_0),
    .io_out_b_0(mesh_1_7_io_out_b_0),
    .io_out_control_0_propagate(mesh_1_7_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_1_7_io_out_control_0_shift),
    .io_in_valid_0(mesh_1_7_io_in_valid_0),
    .io_out_valid_0(mesh_1_7_io_out_valid_0)
  );
  Tile mesh_2_0 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177104.4]
    .clock(mesh_2_0_clock),
    .io_in_a_0(mesh_2_0_io_in_a_0),
    .io_in_b_0(mesh_2_0_io_in_b_0),
    .io_in_d_0(mesh_2_0_io_in_d_0),
    .io_in_control_0_propagate(mesh_2_0_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_2_0_io_in_control_0_shift),
    .io_out_a_0(mesh_2_0_io_out_a_0),
    .io_out_c_0(mesh_2_0_io_out_c_0),
    .io_out_b_0(mesh_2_0_io_out_b_0),
    .io_out_control_0_propagate(mesh_2_0_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_2_0_io_out_control_0_shift),
    .io_in_valid_0(mesh_2_0_io_in_valid_0),
    .io_out_valid_0(mesh_2_0_io_out_valid_0)
  );
  Tile mesh_2_1 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177107.4]
    .clock(mesh_2_1_clock),
    .io_in_a_0(mesh_2_1_io_in_a_0),
    .io_in_b_0(mesh_2_1_io_in_b_0),
    .io_in_d_0(mesh_2_1_io_in_d_0),
    .io_in_control_0_propagate(mesh_2_1_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_2_1_io_in_control_0_shift),
    .io_out_a_0(mesh_2_1_io_out_a_0),
    .io_out_c_0(mesh_2_1_io_out_c_0),
    .io_out_b_0(mesh_2_1_io_out_b_0),
    .io_out_control_0_propagate(mesh_2_1_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_2_1_io_out_control_0_shift),
    .io_in_valid_0(mesh_2_1_io_in_valid_0),
    .io_out_valid_0(mesh_2_1_io_out_valid_0)
  );
  Tile mesh_2_2 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177110.4]
    .clock(mesh_2_2_clock),
    .io_in_a_0(mesh_2_2_io_in_a_0),
    .io_in_b_0(mesh_2_2_io_in_b_0),
    .io_in_d_0(mesh_2_2_io_in_d_0),
    .io_in_control_0_propagate(mesh_2_2_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_2_2_io_in_control_0_shift),
    .io_out_a_0(mesh_2_2_io_out_a_0),
    .io_out_c_0(mesh_2_2_io_out_c_0),
    .io_out_b_0(mesh_2_2_io_out_b_0),
    .io_out_control_0_propagate(mesh_2_2_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_2_2_io_out_control_0_shift),
    .io_in_valid_0(mesh_2_2_io_in_valid_0),
    .io_out_valid_0(mesh_2_2_io_out_valid_0)
  );
  Tile mesh_2_3 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177113.4]
    .clock(mesh_2_3_clock),
    .io_in_a_0(mesh_2_3_io_in_a_0),
    .io_in_b_0(mesh_2_3_io_in_b_0),
    .io_in_d_0(mesh_2_3_io_in_d_0),
    .io_in_control_0_propagate(mesh_2_3_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_2_3_io_in_control_0_shift),
    .io_out_a_0(mesh_2_3_io_out_a_0),
    .io_out_c_0(mesh_2_3_io_out_c_0),
    .io_out_b_0(mesh_2_3_io_out_b_0),
    .io_out_control_0_propagate(mesh_2_3_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_2_3_io_out_control_0_shift),
    .io_in_valid_0(mesh_2_3_io_in_valid_0),
    .io_out_valid_0(mesh_2_3_io_out_valid_0)
  );
  Tile mesh_2_4 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177116.4]
    .clock(mesh_2_4_clock),
    .io_in_a_0(mesh_2_4_io_in_a_0),
    .io_in_b_0(mesh_2_4_io_in_b_0),
    .io_in_d_0(mesh_2_4_io_in_d_0),
    .io_in_control_0_propagate(mesh_2_4_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_2_4_io_in_control_0_shift),
    .io_out_a_0(mesh_2_4_io_out_a_0),
    .io_out_c_0(mesh_2_4_io_out_c_0),
    .io_out_b_0(mesh_2_4_io_out_b_0),
    .io_out_control_0_propagate(mesh_2_4_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_2_4_io_out_control_0_shift),
    .io_in_valid_0(mesh_2_4_io_in_valid_0),
    .io_out_valid_0(mesh_2_4_io_out_valid_0)
  );
  Tile mesh_2_5 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177119.4]
    .clock(mesh_2_5_clock),
    .io_in_a_0(mesh_2_5_io_in_a_0),
    .io_in_b_0(mesh_2_5_io_in_b_0),
    .io_in_d_0(mesh_2_5_io_in_d_0),
    .io_in_control_0_propagate(mesh_2_5_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_2_5_io_in_control_0_shift),
    .io_out_a_0(mesh_2_5_io_out_a_0),
    .io_out_c_0(mesh_2_5_io_out_c_0),
    .io_out_b_0(mesh_2_5_io_out_b_0),
    .io_out_control_0_propagate(mesh_2_5_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_2_5_io_out_control_0_shift),
    .io_in_valid_0(mesh_2_5_io_in_valid_0),
    .io_out_valid_0(mesh_2_5_io_out_valid_0)
  );
  Tile mesh_2_6 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177122.4]
    .clock(mesh_2_6_clock),
    .io_in_a_0(mesh_2_6_io_in_a_0),
    .io_in_b_0(mesh_2_6_io_in_b_0),
    .io_in_d_0(mesh_2_6_io_in_d_0),
    .io_in_control_0_propagate(mesh_2_6_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_2_6_io_in_control_0_shift),
    .io_out_a_0(mesh_2_6_io_out_a_0),
    .io_out_c_0(mesh_2_6_io_out_c_0),
    .io_out_b_0(mesh_2_6_io_out_b_0),
    .io_out_control_0_propagate(mesh_2_6_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_2_6_io_out_control_0_shift),
    .io_in_valid_0(mesh_2_6_io_in_valid_0),
    .io_out_valid_0(mesh_2_6_io_out_valid_0)
  );
  Tile mesh_2_7 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177125.4]
    .clock(mesh_2_7_clock),
    .io_in_a_0(mesh_2_7_io_in_a_0),
    .io_in_b_0(mesh_2_7_io_in_b_0),
    .io_in_d_0(mesh_2_7_io_in_d_0),
    .io_in_control_0_propagate(mesh_2_7_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_2_7_io_in_control_0_shift),
    .io_out_a_0(mesh_2_7_io_out_a_0),
    .io_out_c_0(mesh_2_7_io_out_c_0),
    .io_out_b_0(mesh_2_7_io_out_b_0),
    .io_out_control_0_propagate(mesh_2_7_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_2_7_io_out_control_0_shift),
    .io_in_valid_0(mesh_2_7_io_in_valid_0),
    .io_out_valid_0(mesh_2_7_io_out_valid_0)
  );
  Tile mesh_3_0 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177128.4]
    .clock(mesh_3_0_clock),
    .io_in_a_0(mesh_3_0_io_in_a_0),
    .io_in_b_0(mesh_3_0_io_in_b_0),
    .io_in_d_0(mesh_3_0_io_in_d_0),
    .io_in_control_0_propagate(mesh_3_0_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_3_0_io_in_control_0_shift),
    .io_out_a_0(mesh_3_0_io_out_a_0),
    .io_out_c_0(mesh_3_0_io_out_c_0),
    .io_out_b_0(mesh_3_0_io_out_b_0),
    .io_out_control_0_propagate(mesh_3_0_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_3_0_io_out_control_0_shift),
    .io_in_valid_0(mesh_3_0_io_in_valid_0),
    .io_out_valid_0(mesh_3_0_io_out_valid_0)
  );
  Tile mesh_3_1 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177131.4]
    .clock(mesh_3_1_clock),
    .io_in_a_0(mesh_3_1_io_in_a_0),
    .io_in_b_0(mesh_3_1_io_in_b_0),
    .io_in_d_0(mesh_3_1_io_in_d_0),
    .io_in_control_0_propagate(mesh_3_1_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_3_1_io_in_control_0_shift),
    .io_out_a_0(mesh_3_1_io_out_a_0),
    .io_out_c_0(mesh_3_1_io_out_c_0),
    .io_out_b_0(mesh_3_1_io_out_b_0),
    .io_out_control_0_propagate(mesh_3_1_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_3_1_io_out_control_0_shift),
    .io_in_valid_0(mesh_3_1_io_in_valid_0),
    .io_out_valid_0(mesh_3_1_io_out_valid_0)
  );
  Tile mesh_3_2 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177134.4]
    .clock(mesh_3_2_clock),
    .io_in_a_0(mesh_3_2_io_in_a_0),
    .io_in_b_0(mesh_3_2_io_in_b_0),
    .io_in_d_0(mesh_3_2_io_in_d_0),
    .io_in_control_0_propagate(mesh_3_2_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_3_2_io_in_control_0_shift),
    .io_out_a_0(mesh_3_2_io_out_a_0),
    .io_out_c_0(mesh_3_2_io_out_c_0),
    .io_out_b_0(mesh_3_2_io_out_b_0),
    .io_out_control_0_propagate(mesh_3_2_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_3_2_io_out_control_0_shift),
    .io_in_valid_0(mesh_3_2_io_in_valid_0),
    .io_out_valid_0(mesh_3_2_io_out_valid_0)
  );
  Tile mesh_3_3 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177137.4]
    .clock(mesh_3_3_clock),
    .io_in_a_0(mesh_3_3_io_in_a_0),
    .io_in_b_0(mesh_3_3_io_in_b_0),
    .io_in_d_0(mesh_3_3_io_in_d_0),
    .io_in_control_0_propagate(mesh_3_3_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_3_3_io_in_control_0_shift),
    .io_out_a_0(mesh_3_3_io_out_a_0),
    .io_out_c_0(mesh_3_3_io_out_c_0),
    .io_out_b_0(mesh_3_3_io_out_b_0),
    .io_out_control_0_propagate(mesh_3_3_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_3_3_io_out_control_0_shift),
    .io_in_valid_0(mesh_3_3_io_in_valid_0),
    .io_out_valid_0(mesh_3_3_io_out_valid_0)
  );
  Tile mesh_3_4 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177140.4]
    .clock(mesh_3_4_clock),
    .io_in_a_0(mesh_3_4_io_in_a_0),
    .io_in_b_0(mesh_3_4_io_in_b_0),
    .io_in_d_0(mesh_3_4_io_in_d_0),
    .io_in_control_0_propagate(mesh_3_4_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_3_4_io_in_control_0_shift),
    .io_out_a_0(mesh_3_4_io_out_a_0),
    .io_out_c_0(mesh_3_4_io_out_c_0),
    .io_out_b_0(mesh_3_4_io_out_b_0),
    .io_out_control_0_propagate(mesh_3_4_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_3_4_io_out_control_0_shift),
    .io_in_valid_0(mesh_3_4_io_in_valid_0),
    .io_out_valid_0(mesh_3_4_io_out_valid_0)
  );
  Tile mesh_3_5 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177143.4]
    .clock(mesh_3_5_clock),
    .io_in_a_0(mesh_3_5_io_in_a_0),
    .io_in_b_0(mesh_3_5_io_in_b_0),
    .io_in_d_0(mesh_3_5_io_in_d_0),
    .io_in_control_0_propagate(mesh_3_5_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_3_5_io_in_control_0_shift),
    .io_out_a_0(mesh_3_5_io_out_a_0),
    .io_out_c_0(mesh_3_5_io_out_c_0),
    .io_out_b_0(mesh_3_5_io_out_b_0),
    .io_out_control_0_propagate(mesh_3_5_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_3_5_io_out_control_0_shift),
    .io_in_valid_0(mesh_3_5_io_in_valid_0),
    .io_out_valid_0(mesh_3_5_io_out_valid_0)
  );
  Tile mesh_3_6 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177146.4]
    .clock(mesh_3_6_clock),
    .io_in_a_0(mesh_3_6_io_in_a_0),
    .io_in_b_0(mesh_3_6_io_in_b_0),
    .io_in_d_0(mesh_3_6_io_in_d_0),
    .io_in_control_0_propagate(mesh_3_6_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_3_6_io_in_control_0_shift),
    .io_out_a_0(mesh_3_6_io_out_a_0),
    .io_out_c_0(mesh_3_6_io_out_c_0),
    .io_out_b_0(mesh_3_6_io_out_b_0),
    .io_out_control_0_propagate(mesh_3_6_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_3_6_io_out_control_0_shift),
    .io_in_valid_0(mesh_3_6_io_in_valid_0),
    .io_out_valid_0(mesh_3_6_io_out_valid_0)
  );
  Tile mesh_3_7 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177149.4]
    .clock(mesh_3_7_clock),
    .io_in_a_0(mesh_3_7_io_in_a_0),
    .io_in_b_0(mesh_3_7_io_in_b_0),
    .io_in_d_0(mesh_3_7_io_in_d_0),
    .io_in_control_0_propagate(mesh_3_7_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_3_7_io_in_control_0_shift),
    .io_out_a_0(mesh_3_7_io_out_a_0),
    .io_out_c_0(mesh_3_7_io_out_c_0),
    .io_out_b_0(mesh_3_7_io_out_b_0),
    .io_out_control_0_propagate(mesh_3_7_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_3_7_io_out_control_0_shift),
    .io_in_valid_0(mesh_3_7_io_in_valid_0),
    .io_out_valid_0(mesh_3_7_io_out_valid_0)
  );
  Tile mesh_4_0 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177152.4]
    .clock(mesh_4_0_clock),
    .io_in_a_0(mesh_4_0_io_in_a_0),
    .io_in_b_0(mesh_4_0_io_in_b_0),
    .io_in_d_0(mesh_4_0_io_in_d_0),
    .io_in_control_0_propagate(mesh_4_0_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_4_0_io_in_control_0_shift),
    .io_out_a_0(mesh_4_0_io_out_a_0),
    .io_out_c_0(mesh_4_0_io_out_c_0),
    .io_out_b_0(mesh_4_0_io_out_b_0),
    .io_out_control_0_propagate(mesh_4_0_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_4_0_io_out_control_0_shift),
    .io_in_valid_0(mesh_4_0_io_in_valid_0),
    .io_out_valid_0(mesh_4_0_io_out_valid_0)
  );
  Tile mesh_4_1 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177155.4]
    .clock(mesh_4_1_clock),
    .io_in_a_0(mesh_4_1_io_in_a_0),
    .io_in_b_0(mesh_4_1_io_in_b_0),
    .io_in_d_0(mesh_4_1_io_in_d_0),
    .io_in_control_0_propagate(mesh_4_1_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_4_1_io_in_control_0_shift),
    .io_out_a_0(mesh_4_1_io_out_a_0),
    .io_out_c_0(mesh_4_1_io_out_c_0),
    .io_out_b_0(mesh_4_1_io_out_b_0),
    .io_out_control_0_propagate(mesh_4_1_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_4_1_io_out_control_0_shift),
    .io_in_valid_0(mesh_4_1_io_in_valid_0),
    .io_out_valid_0(mesh_4_1_io_out_valid_0)
  );
  Tile mesh_4_2 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177158.4]
    .clock(mesh_4_2_clock),
    .io_in_a_0(mesh_4_2_io_in_a_0),
    .io_in_b_0(mesh_4_2_io_in_b_0),
    .io_in_d_0(mesh_4_2_io_in_d_0),
    .io_in_control_0_propagate(mesh_4_2_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_4_2_io_in_control_0_shift),
    .io_out_a_0(mesh_4_2_io_out_a_0),
    .io_out_c_0(mesh_4_2_io_out_c_0),
    .io_out_b_0(mesh_4_2_io_out_b_0),
    .io_out_control_0_propagate(mesh_4_2_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_4_2_io_out_control_0_shift),
    .io_in_valid_0(mesh_4_2_io_in_valid_0),
    .io_out_valid_0(mesh_4_2_io_out_valid_0)
  );
  Tile mesh_4_3 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177161.4]
    .clock(mesh_4_3_clock),
    .io_in_a_0(mesh_4_3_io_in_a_0),
    .io_in_b_0(mesh_4_3_io_in_b_0),
    .io_in_d_0(mesh_4_3_io_in_d_0),
    .io_in_control_0_propagate(mesh_4_3_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_4_3_io_in_control_0_shift),
    .io_out_a_0(mesh_4_3_io_out_a_0),
    .io_out_c_0(mesh_4_3_io_out_c_0),
    .io_out_b_0(mesh_4_3_io_out_b_0),
    .io_out_control_0_propagate(mesh_4_3_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_4_3_io_out_control_0_shift),
    .io_in_valid_0(mesh_4_3_io_in_valid_0),
    .io_out_valid_0(mesh_4_3_io_out_valid_0)
  );
  Tile mesh_4_4 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177164.4]
    .clock(mesh_4_4_clock),
    .io_in_a_0(mesh_4_4_io_in_a_0),
    .io_in_b_0(mesh_4_4_io_in_b_0),
    .io_in_d_0(mesh_4_4_io_in_d_0),
    .io_in_control_0_propagate(mesh_4_4_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_4_4_io_in_control_0_shift),
    .io_out_a_0(mesh_4_4_io_out_a_0),
    .io_out_c_0(mesh_4_4_io_out_c_0),
    .io_out_b_0(mesh_4_4_io_out_b_0),
    .io_out_control_0_propagate(mesh_4_4_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_4_4_io_out_control_0_shift),
    .io_in_valid_0(mesh_4_4_io_in_valid_0),
    .io_out_valid_0(mesh_4_4_io_out_valid_0)
  );
  Tile mesh_4_5 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177167.4]
    .clock(mesh_4_5_clock),
    .io_in_a_0(mesh_4_5_io_in_a_0),
    .io_in_b_0(mesh_4_5_io_in_b_0),
    .io_in_d_0(mesh_4_5_io_in_d_0),
    .io_in_control_0_propagate(mesh_4_5_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_4_5_io_in_control_0_shift),
    .io_out_a_0(mesh_4_5_io_out_a_0),
    .io_out_c_0(mesh_4_5_io_out_c_0),
    .io_out_b_0(mesh_4_5_io_out_b_0),
    .io_out_control_0_propagate(mesh_4_5_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_4_5_io_out_control_0_shift),
    .io_in_valid_0(mesh_4_5_io_in_valid_0),
    .io_out_valid_0(mesh_4_5_io_out_valid_0)
  );
  Tile mesh_4_6 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177170.4]
    .clock(mesh_4_6_clock),
    .io_in_a_0(mesh_4_6_io_in_a_0),
    .io_in_b_0(mesh_4_6_io_in_b_0),
    .io_in_d_0(mesh_4_6_io_in_d_0),
    .io_in_control_0_propagate(mesh_4_6_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_4_6_io_in_control_0_shift),
    .io_out_a_0(mesh_4_6_io_out_a_0),
    .io_out_c_0(mesh_4_6_io_out_c_0),
    .io_out_b_0(mesh_4_6_io_out_b_0),
    .io_out_control_0_propagate(mesh_4_6_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_4_6_io_out_control_0_shift),
    .io_in_valid_0(mesh_4_6_io_in_valid_0),
    .io_out_valid_0(mesh_4_6_io_out_valid_0)
  );
  Tile mesh_4_7 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177173.4]
    .clock(mesh_4_7_clock),
    .io_in_a_0(mesh_4_7_io_in_a_0),
    .io_in_b_0(mesh_4_7_io_in_b_0),
    .io_in_d_0(mesh_4_7_io_in_d_0),
    .io_in_control_0_propagate(mesh_4_7_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_4_7_io_in_control_0_shift),
    .io_out_a_0(mesh_4_7_io_out_a_0),
    .io_out_c_0(mesh_4_7_io_out_c_0),
    .io_out_b_0(mesh_4_7_io_out_b_0),
    .io_out_control_0_propagate(mesh_4_7_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_4_7_io_out_control_0_shift),
    .io_in_valid_0(mesh_4_7_io_in_valid_0),
    .io_out_valid_0(mesh_4_7_io_out_valid_0)
  );
  Tile mesh_5_0 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177176.4]
    .clock(mesh_5_0_clock),
    .io_in_a_0(mesh_5_0_io_in_a_0),
    .io_in_b_0(mesh_5_0_io_in_b_0),
    .io_in_d_0(mesh_5_0_io_in_d_0),
    .io_in_control_0_propagate(mesh_5_0_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_5_0_io_in_control_0_shift),
    .io_out_a_0(mesh_5_0_io_out_a_0),
    .io_out_c_0(mesh_5_0_io_out_c_0),
    .io_out_b_0(mesh_5_0_io_out_b_0),
    .io_out_control_0_propagate(mesh_5_0_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_5_0_io_out_control_0_shift),
    .io_in_valid_0(mesh_5_0_io_in_valid_0),
    .io_out_valid_0(mesh_5_0_io_out_valid_0)
  );
  Tile mesh_5_1 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177179.4]
    .clock(mesh_5_1_clock),
    .io_in_a_0(mesh_5_1_io_in_a_0),
    .io_in_b_0(mesh_5_1_io_in_b_0),
    .io_in_d_0(mesh_5_1_io_in_d_0),
    .io_in_control_0_propagate(mesh_5_1_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_5_1_io_in_control_0_shift),
    .io_out_a_0(mesh_5_1_io_out_a_0),
    .io_out_c_0(mesh_5_1_io_out_c_0),
    .io_out_b_0(mesh_5_1_io_out_b_0),
    .io_out_control_0_propagate(mesh_5_1_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_5_1_io_out_control_0_shift),
    .io_in_valid_0(mesh_5_1_io_in_valid_0),
    .io_out_valid_0(mesh_5_1_io_out_valid_0)
  );
  Tile mesh_5_2 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177182.4]
    .clock(mesh_5_2_clock),
    .io_in_a_0(mesh_5_2_io_in_a_0),
    .io_in_b_0(mesh_5_2_io_in_b_0),
    .io_in_d_0(mesh_5_2_io_in_d_0),
    .io_in_control_0_propagate(mesh_5_2_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_5_2_io_in_control_0_shift),
    .io_out_a_0(mesh_5_2_io_out_a_0),
    .io_out_c_0(mesh_5_2_io_out_c_0),
    .io_out_b_0(mesh_5_2_io_out_b_0),
    .io_out_control_0_propagate(mesh_5_2_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_5_2_io_out_control_0_shift),
    .io_in_valid_0(mesh_5_2_io_in_valid_0),
    .io_out_valid_0(mesh_5_2_io_out_valid_0)
  );
  Tile mesh_5_3 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177185.4]
    .clock(mesh_5_3_clock),
    .io_in_a_0(mesh_5_3_io_in_a_0),
    .io_in_b_0(mesh_5_3_io_in_b_0),
    .io_in_d_0(mesh_5_3_io_in_d_0),
    .io_in_control_0_propagate(mesh_5_3_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_5_3_io_in_control_0_shift),
    .io_out_a_0(mesh_5_3_io_out_a_0),
    .io_out_c_0(mesh_5_3_io_out_c_0),
    .io_out_b_0(mesh_5_3_io_out_b_0),
    .io_out_control_0_propagate(mesh_5_3_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_5_3_io_out_control_0_shift),
    .io_in_valid_0(mesh_5_3_io_in_valid_0),
    .io_out_valid_0(mesh_5_3_io_out_valid_0)
  );
  Tile mesh_5_4 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177188.4]
    .clock(mesh_5_4_clock),
    .io_in_a_0(mesh_5_4_io_in_a_0),
    .io_in_b_0(mesh_5_4_io_in_b_0),
    .io_in_d_0(mesh_5_4_io_in_d_0),
    .io_in_control_0_propagate(mesh_5_4_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_5_4_io_in_control_0_shift),
    .io_out_a_0(mesh_5_4_io_out_a_0),
    .io_out_c_0(mesh_5_4_io_out_c_0),
    .io_out_b_0(mesh_5_4_io_out_b_0),
    .io_out_control_0_propagate(mesh_5_4_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_5_4_io_out_control_0_shift),
    .io_in_valid_0(mesh_5_4_io_in_valid_0),
    .io_out_valid_0(mesh_5_4_io_out_valid_0)
  );
  Tile mesh_5_5 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177191.4]
    .clock(mesh_5_5_clock),
    .io_in_a_0(mesh_5_5_io_in_a_0),
    .io_in_b_0(mesh_5_5_io_in_b_0),
    .io_in_d_0(mesh_5_5_io_in_d_0),
    .io_in_control_0_propagate(mesh_5_5_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_5_5_io_in_control_0_shift),
    .io_out_a_0(mesh_5_5_io_out_a_0),
    .io_out_c_0(mesh_5_5_io_out_c_0),
    .io_out_b_0(mesh_5_5_io_out_b_0),
    .io_out_control_0_propagate(mesh_5_5_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_5_5_io_out_control_0_shift),
    .io_in_valid_0(mesh_5_5_io_in_valid_0),
    .io_out_valid_0(mesh_5_5_io_out_valid_0)
  );
  Tile mesh_5_6 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177194.4]
    .clock(mesh_5_6_clock),
    .io_in_a_0(mesh_5_6_io_in_a_0),
    .io_in_b_0(mesh_5_6_io_in_b_0),
    .io_in_d_0(mesh_5_6_io_in_d_0),
    .io_in_control_0_propagate(mesh_5_6_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_5_6_io_in_control_0_shift),
    .io_out_a_0(mesh_5_6_io_out_a_0),
    .io_out_c_0(mesh_5_6_io_out_c_0),
    .io_out_b_0(mesh_5_6_io_out_b_0),
    .io_out_control_0_propagate(mesh_5_6_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_5_6_io_out_control_0_shift),
    .io_in_valid_0(mesh_5_6_io_in_valid_0),
    .io_out_valid_0(mesh_5_6_io_out_valid_0)
  );
  Tile mesh_5_7 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177197.4]
    .clock(mesh_5_7_clock),
    .io_in_a_0(mesh_5_7_io_in_a_0),
    .io_in_b_0(mesh_5_7_io_in_b_0),
    .io_in_d_0(mesh_5_7_io_in_d_0),
    .io_in_control_0_propagate(mesh_5_7_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_5_7_io_in_control_0_shift),
    .io_out_a_0(mesh_5_7_io_out_a_0),
    .io_out_c_0(mesh_5_7_io_out_c_0),
    .io_out_b_0(mesh_5_7_io_out_b_0),
    .io_out_control_0_propagate(mesh_5_7_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_5_7_io_out_control_0_shift),
    .io_in_valid_0(mesh_5_7_io_in_valid_0),
    .io_out_valid_0(mesh_5_7_io_out_valid_0)
  );
  Tile mesh_6_0 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177200.4]
    .clock(mesh_6_0_clock),
    .io_in_a_0(mesh_6_0_io_in_a_0),
    .io_in_b_0(mesh_6_0_io_in_b_0),
    .io_in_d_0(mesh_6_0_io_in_d_0),
    .io_in_control_0_propagate(mesh_6_0_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_6_0_io_in_control_0_shift),
    .io_out_a_0(mesh_6_0_io_out_a_0),
    .io_out_c_0(mesh_6_0_io_out_c_0),
    .io_out_b_0(mesh_6_0_io_out_b_0),
    .io_out_control_0_propagate(mesh_6_0_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_6_0_io_out_control_0_shift),
    .io_in_valid_0(mesh_6_0_io_in_valid_0),
    .io_out_valid_0(mesh_6_0_io_out_valid_0)
  );
  Tile mesh_6_1 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177203.4]
    .clock(mesh_6_1_clock),
    .io_in_a_0(mesh_6_1_io_in_a_0),
    .io_in_b_0(mesh_6_1_io_in_b_0),
    .io_in_d_0(mesh_6_1_io_in_d_0),
    .io_in_control_0_propagate(mesh_6_1_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_6_1_io_in_control_0_shift),
    .io_out_a_0(mesh_6_1_io_out_a_0),
    .io_out_c_0(mesh_6_1_io_out_c_0),
    .io_out_b_0(mesh_6_1_io_out_b_0),
    .io_out_control_0_propagate(mesh_6_1_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_6_1_io_out_control_0_shift),
    .io_in_valid_0(mesh_6_1_io_in_valid_0),
    .io_out_valid_0(mesh_6_1_io_out_valid_0)
  );
  Tile mesh_6_2 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177206.4]
    .clock(mesh_6_2_clock),
    .io_in_a_0(mesh_6_2_io_in_a_0),
    .io_in_b_0(mesh_6_2_io_in_b_0),
    .io_in_d_0(mesh_6_2_io_in_d_0),
    .io_in_control_0_propagate(mesh_6_2_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_6_2_io_in_control_0_shift),
    .io_out_a_0(mesh_6_2_io_out_a_0),
    .io_out_c_0(mesh_6_2_io_out_c_0),
    .io_out_b_0(mesh_6_2_io_out_b_0),
    .io_out_control_0_propagate(mesh_6_2_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_6_2_io_out_control_0_shift),
    .io_in_valid_0(mesh_6_2_io_in_valid_0),
    .io_out_valid_0(mesh_6_2_io_out_valid_0)
  );
  Tile mesh_6_3 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177209.4]
    .clock(mesh_6_3_clock),
    .io_in_a_0(mesh_6_3_io_in_a_0),
    .io_in_b_0(mesh_6_3_io_in_b_0),
    .io_in_d_0(mesh_6_3_io_in_d_0),
    .io_in_control_0_propagate(mesh_6_3_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_6_3_io_in_control_0_shift),
    .io_out_a_0(mesh_6_3_io_out_a_0),
    .io_out_c_0(mesh_6_3_io_out_c_0),
    .io_out_b_0(mesh_6_3_io_out_b_0),
    .io_out_control_0_propagate(mesh_6_3_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_6_3_io_out_control_0_shift),
    .io_in_valid_0(mesh_6_3_io_in_valid_0),
    .io_out_valid_0(mesh_6_3_io_out_valid_0)
  );
  Tile mesh_6_4 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177212.4]
    .clock(mesh_6_4_clock),
    .io_in_a_0(mesh_6_4_io_in_a_0),
    .io_in_b_0(mesh_6_4_io_in_b_0),
    .io_in_d_0(mesh_6_4_io_in_d_0),
    .io_in_control_0_propagate(mesh_6_4_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_6_4_io_in_control_0_shift),
    .io_out_a_0(mesh_6_4_io_out_a_0),
    .io_out_c_0(mesh_6_4_io_out_c_0),
    .io_out_b_0(mesh_6_4_io_out_b_0),
    .io_out_control_0_propagate(mesh_6_4_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_6_4_io_out_control_0_shift),
    .io_in_valid_0(mesh_6_4_io_in_valid_0),
    .io_out_valid_0(mesh_6_4_io_out_valid_0)
  );
  Tile mesh_6_5 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177215.4]
    .clock(mesh_6_5_clock),
    .io_in_a_0(mesh_6_5_io_in_a_0),
    .io_in_b_0(mesh_6_5_io_in_b_0),
    .io_in_d_0(mesh_6_5_io_in_d_0),
    .io_in_control_0_propagate(mesh_6_5_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_6_5_io_in_control_0_shift),
    .io_out_a_0(mesh_6_5_io_out_a_0),
    .io_out_c_0(mesh_6_5_io_out_c_0),
    .io_out_b_0(mesh_6_5_io_out_b_0),
    .io_out_control_0_propagate(mesh_6_5_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_6_5_io_out_control_0_shift),
    .io_in_valid_0(mesh_6_5_io_in_valid_0),
    .io_out_valid_0(mesh_6_5_io_out_valid_0)
  );
  Tile mesh_6_6 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177218.4]
    .clock(mesh_6_6_clock),
    .io_in_a_0(mesh_6_6_io_in_a_0),
    .io_in_b_0(mesh_6_6_io_in_b_0),
    .io_in_d_0(mesh_6_6_io_in_d_0),
    .io_in_control_0_propagate(mesh_6_6_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_6_6_io_in_control_0_shift),
    .io_out_a_0(mesh_6_6_io_out_a_0),
    .io_out_c_0(mesh_6_6_io_out_c_0),
    .io_out_b_0(mesh_6_6_io_out_b_0),
    .io_out_control_0_propagate(mesh_6_6_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_6_6_io_out_control_0_shift),
    .io_in_valid_0(mesh_6_6_io_in_valid_0),
    .io_out_valid_0(mesh_6_6_io_out_valid_0)
  );
  Tile mesh_6_7 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177221.4]
    .clock(mesh_6_7_clock),
    .io_in_a_0(mesh_6_7_io_in_a_0),
    .io_in_b_0(mesh_6_7_io_in_b_0),
    .io_in_d_0(mesh_6_7_io_in_d_0),
    .io_in_control_0_propagate(mesh_6_7_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_6_7_io_in_control_0_shift),
    .io_out_a_0(mesh_6_7_io_out_a_0),
    .io_out_c_0(mesh_6_7_io_out_c_0),
    .io_out_b_0(mesh_6_7_io_out_b_0),
    .io_out_control_0_propagate(mesh_6_7_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_6_7_io_out_control_0_shift),
    .io_in_valid_0(mesh_6_7_io_in_valid_0),
    .io_out_valid_0(mesh_6_7_io_out_valid_0)
  );
  Tile mesh_7_0 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177224.4]
    .clock(mesh_7_0_clock),
    .io_in_a_0(mesh_7_0_io_in_a_0),
    .io_in_b_0(mesh_7_0_io_in_b_0),
    .io_in_d_0(mesh_7_0_io_in_d_0),
    .io_in_control_0_propagate(mesh_7_0_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_7_0_io_in_control_0_shift),
    .io_out_a_0(mesh_7_0_io_out_a_0),
    .io_out_c_0(mesh_7_0_io_out_c_0),
    .io_out_b_0(mesh_7_0_io_out_b_0),
    .io_out_control_0_propagate(mesh_7_0_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_7_0_io_out_control_0_shift),
    .io_in_valid_0(mesh_7_0_io_in_valid_0),
    .io_out_valid_0(mesh_7_0_io_out_valid_0)
  );
  Tile mesh_7_1 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177227.4]
    .clock(mesh_7_1_clock),
    .io_in_a_0(mesh_7_1_io_in_a_0),
    .io_in_b_0(mesh_7_1_io_in_b_0),
    .io_in_d_0(mesh_7_1_io_in_d_0),
    .io_in_control_0_propagate(mesh_7_1_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_7_1_io_in_control_0_shift),
    .io_out_a_0(mesh_7_1_io_out_a_0),
    .io_out_c_0(mesh_7_1_io_out_c_0),
    .io_out_b_0(mesh_7_1_io_out_b_0),
    .io_out_control_0_propagate(mesh_7_1_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_7_1_io_out_control_0_shift),
    .io_in_valid_0(mesh_7_1_io_in_valid_0),
    .io_out_valid_0(mesh_7_1_io_out_valid_0)
  );
  Tile mesh_7_2 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177230.4]
    .clock(mesh_7_2_clock),
    .io_in_a_0(mesh_7_2_io_in_a_0),
    .io_in_b_0(mesh_7_2_io_in_b_0),
    .io_in_d_0(mesh_7_2_io_in_d_0),
    .io_in_control_0_propagate(mesh_7_2_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_7_2_io_in_control_0_shift),
    .io_out_a_0(mesh_7_2_io_out_a_0),
    .io_out_c_0(mesh_7_2_io_out_c_0),
    .io_out_b_0(mesh_7_2_io_out_b_0),
    .io_out_control_0_propagate(mesh_7_2_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_7_2_io_out_control_0_shift),
    .io_in_valid_0(mesh_7_2_io_in_valid_0),
    .io_out_valid_0(mesh_7_2_io_out_valid_0)
  );
  Tile mesh_7_3 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177233.4]
    .clock(mesh_7_3_clock),
    .io_in_a_0(mesh_7_3_io_in_a_0),
    .io_in_b_0(mesh_7_3_io_in_b_0),
    .io_in_d_0(mesh_7_3_io_in_d_0),
    .io_in_control_0_propagate(mesh_7_3_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_7_3_io_in_control_0_shift),
    .io_out_a_0(mesh_7_3_io_out_a_0),
    .io_out_c_0(mesh_7_3_io_out_c_0),
    .io_out_b_0(mesh_7_3_io_out_b_0),
    .io_out_control_0_propagate(mesh_7_3_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_7_3_io_out_control_0_shift),
    .io_in_valid_0(mesh_7_3_io_in_valid_0),
    .io_out_valid_0(mesh_7_3_io_out_valid_0)
  );
  Tile mesh_7_4 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177236.4]
    .clock(mesh_7_4_clock),
    .io_in_a_0(mesh_7_4_io_in_a_0),
    .io_in_b_0(mesh_7_4_io_in_b_0),
    .io_in_d_0(mesh_7_4_io_in_d_0),
    .io_in_control_0_propagate(mesh_7_4_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_7_4_io_in_control_0_shift),
    .io_out_a_0(mesh_7_4_io_out_a_0),
    .io_out_c_0(mesh_7_4_io_out_c_0),
    .io_out_b_0(mesh_7_4_io_out_b_0),
    .io_out_control_0_propagate(mesh_7_4_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_7_4_io_out_control_0_shift),
    .io_in_valid_0(mesh_7_4_io_in_valid_0),
    .io_out_valid_0(mesh_7_4_io_out_valid_0)
  );
  Tile mesh_7_5 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177239.4]
    .clock(mesh_7_5_clock),
    .io_in_a_0(mesh_7_5_io_in_a_0),
    .io_in_b_0(mesh_7_5_io_in_b_0),
    .io_in_d_0(mesh_7_5_io_in_d_0),
    .io_in_control_0_propagate(mesh_7_5_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_7_5_io_in_control_0_shift),
    .io_out_a_0(mesh_7_5_io_out_a_0),
    .io_out_c_0(mesh_7_5_io_out_c_0),
    .io_out_b_0(mesh_7_5_io_out_b_0),
    .io_out_control_0_propagate(mesh_7_5_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_7_5_io_out_control_0_shift),
    .io_in_valid_0(mesh_7_5_io_in_valid_0),
    .io_out_valid_0(mesh_7_5_io_out_valid_0)
  );
  Tile mesh_7_6 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177242.4]
    .clock(mesh_7_6_clock),
    .io_in_a_0(mesh_7_6_io_in_a_0),
    .io_in_b_0(mesh_7_6_io_in_b_0),
    .io_in_d_0(mesh_7_6_io_in_d_0),
    .io_in_control_0_propagate(mesh_7_6_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_7_6_io_in_control_0_shift),
    .io_out_a_0(mesh_7_6_io_out_a_0),
    .io_out_c_0(mesh_7_6_io_out_c_0),
    .io_out_b_0(mesh_7_6_io_out_b_0),
    .io_out_control_0_propagate(mesh_7_6_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_7_6_io_out_control_0_shift),
    .io_in_valid_0(mesh_7_6_io_in_valid_0),
    .io_out_valid_0(mesh_7_6_io_out_valid_0)
  );
  Tile mesh_7_7 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig.fir@177245.4]
    .clock(mesh_7_7_clock),
    .io_in_a_0(mesh_7_7_io_in_a_0),
    .io_in_b_0(mesh_7_7_io_in_b_0),
    .io_in_d_0(mesh_7_7_io_in_d_0),
    .io_in_control_0_propagate(mesh_7_7_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_7_7_io_in_control_0_shift),
    .io_out_a_0(mesh_7_7_io_out_a_0),
    .io_out_c_0(mesh_7_7_io_out_c_0),
    .io_out_b_0(mesh_7_7_io_out_b_0),
    .io_out_control_0_propagate(mesh_7_7_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_7_7_io_out_control_0_shift),
    .io_in_valid_0(mesh_7_7_io_in_valid_0),
    .io_out_valid_0(mesh_7_7_io_out_valid_0)
  );
  assign io_out_c_0_0 = mesh_7_0_io_out_b_0; // @[Mesh.scala 85:7:example.TestHarness.GemminiSocTest1RocketConfig.fir@179376.4]
  assign io_out_c_1_0 = mesh_7_1_io_out_b_0; // @[Mesh.scala 85:7:example.TestHarness.GemminiSocTest1RocketConfig.fir@179379.4]
  assign io_out_c_2_0 = mesh_7_2_io_out_b_0; // @[Mesh.scala 85:7:example.TestHarness.GemminiSocTest1RocketConfig.fir@179382.4]
  assign io_out_c_3_0 = mesh_7_3_io_out_b_0; // @[Mesh.scala 85:7:example.TestHarness.GemminiSocTest1RocketConfig.fir@179385.4]
  assign io_out_c_4_0 = mesh_7_4_io_out_b_0; // @[Mesh.scala 85:7:example.TestHarness.GemminiSocTest1RocketConfig.fir@179388.4]
  assign io_out_c_5_0 = mesh_7_5_io_out_b_0; // @[Mesh.scala 85:7:example.TestHarness.GemminiSocTest1RocketConfig.fir@179391.4]
  assign io_out_c_6_0 = mesh_7_6_io_out_b_0; // @[Mesh.scala 85:7:example.TestHarness.GemminiSocTest1RocketConfig.fir@179394.4]
  assign io_out_c_7_0 = mesh_7_7_io_out_b_0; // @[Mesh.scala 85:7:example.TestHarness.GemminiSocTest1RocketConfig.fir@179397.4]
  assign io_out_b_0_0 = mesh_7_0_io_out_c_0; // @[Mesh.scala 86:7:example.TestHarness.GemminiSocTest1RocketConfig.fir@179377.4]
  assign io_out_b_1_0 = mesh_7_1_io_out_c_0; // @[Mesh.scala 86:7:example.TestHarness.GemminiSocTest1RocketConfig.fir@179380.4]
  assign io_out_b_2_0 = mesh_7_2_io_out_c_0; // @[Mesh.scala 86:7:example.TestHarness.GemminiSocTest1RocketConfig.fir@179383.4]
  assign io_out_b_3_0 = mesh_7_3_io_out_c_0; // @[Mesh.scala 86:7:example.TestHarness.GemminiSocTest1RocketConfig.fir@179386.4]
  assign io_out_b_4_0 = mesh_7_4_io_out_c_0; // @[Mesh.scala 86:7:example.TestHarness.GemminiSocTest1RocketConfig.fir@179389.4]
  assign io_out_b_5_0 = mesh_7_5_io_out_c_0; // @[Mesh.scala 86:7:example.TestHarness.GemminiSocTest1RocketConfig.fir@179392.4]
  assign io_out_b_6_0 = mesh_7_6_io_out_c_0; // @[Mesh.scala 86:7:example.TestHarness.GemminiSocTest1RocketConfig.fir@179395.4]
  assign io_out_b_7_0 = mesh_7_7_io_out_c_0; // @[Mesh.scala 86:7:example.TestHarness.GemminiSocTest1RocketConfig.fir@179398.4]
  assign io_out_valid_0_0 = mesh_7_0_io_out_valid_0; // @[Mesh.scala 87:7:example.TestHarness.GemminiSocTest1RocketConfig.fir@179378.4]
  assign mesh_0_0_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177057.4]
  assign mesh_0_0_io_in_a_0 = _T_1_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177252.4]
  assign mesh_0_0_io_in_b_0 = {{11{_T_74_0[7]}},_T_74_0}; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177464.4]
  assign mesh_0_0_io_in_d_0 = {{11{_T_154_0[7]}},_T_154_0}; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177816.4]
  assign mesh_0_0_io_in_control_0_propagate = _T_236; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178180.4]
  assign mesh_0_0_io_in_control_0_shift = _T_234; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178170.4]
  assign mesh_0_0_io_in_valid_0 = _T_441_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179172.4]
  assign mesh_0_1_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177060.4]
  assign mesh_0_1_io_in_a_0 = _T_2_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177255.4]
  assign mesh_0_1_io_in_b_0 = {{11{_T_84_0[7]}},_T_84_0}; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177508.4]
  assign mesh_0_1_io_in_d_0 = {{11{_T_164_0[7]}},_T_164_0}; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177860.4]
  assign mesh_0_1_io_in_control_0_propagate = _T_262; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178306.4]
  assign mesh_0_1_io_in_control_0_shift = _T_260; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178296.4]
  assign mesh_0_1_io_in_valid_0 = _T_450_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179198.4]
  assign mesh_0_2_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177063.4]
  assign mesh_0_2_io_in_a_0 = _T_3_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177258.4]
  assign mesh_0_2_io_in_b_0 = {{11{_T_94_0[7]}},_T_94_0}; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177552.4]
  assign mesh_0_2_io_in_d_0 = {{11{_T_174_0[7]}},_T_174_0}; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177904.4]
  assign mesh_0_2_io_in_control_0_propagate = _T_288; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178432.4]
  assign mesh_0_2_io_in_control_0_shift = _T_286; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178422.4]
  assign mesh_0_2_io_in_valid_0 = _T_459_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179224.4]
  assign mesh_0_3_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177066.4]
  assign mesh_0_3_io_in_a_0 = _T_4_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177261.4]
  assign mesh_0_3_io_in_b_0 = {{11{_T_104_0[7]}},_T_104_0}; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177596.4]
  assign mesh_0_3_io_in_d_0 = {{11{_T_184_0[7]}},_T_184_0}; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177948.4]
  assign mesh_0_3_io_in_control_0_propagate = _T_314; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178558.4]
  assign mesh_0_3_io_in_control_0_shift = _T_312; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178548.4]
  assign mesh_0_3_io_in_valid_0 = _T_468_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179250.4]
  assign mesh_0_4_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177069.4]
  assign mesh_0_4_io_in_a_0 = _T_5_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177264.4]
  assign mesh_0_4_io_in_b_0 = {{11{_T_114_0[7]}},_T_114_0}; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177640.4]
  assign mesh_0_4_io_in_d_0 = {{11{_T_194_0[7]}},_T_194_0}; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177992.4]
  assign mesh_0_4_io_in_control_0_propagate = _T_340; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178684.4]
  assign mesh_0_4_io_in_control_0_shift = _T_338; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178674.4]
  assign mesh_0_4_io_in_valid_0 = _T_477_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179276.4]
  assign mesh_0_5_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177072.4]
  assign mesh_0_5_io_in_a_0 = _T_6_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177267.4]
  assign mesh_0_5_io_in_b_0 = {{11{_T_124_0[7]}},_T_124_0}; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177684.4]
  assign mesh_0_5_io_in_d_0 = {{11{_T_204_0[7]}},_T_204_0}; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@178036.4]
  assign mesh_0_5_io_in_control_0_propagate = _T_366; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178810.4]
  assign mesh_0_5_io_in_control_0_shift = _T_364; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178800.4]
  assign mesh_0_5_io_in_valid_0 = _T_486_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179302.4]
  assign mesh_0_6_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177075.4]
  assign mesh_0_6_io_in_a_0 = _T_7_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177270.4]
  assign mesh_0_6_io_in_b_0 = {{11{_T_134_0[7]}},_T_134_0}; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177728.4]
  assign mesh_0_6_io_in_d_0 = {{11{_T_214_0[7]}},_T_214_0}; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@178080.4]
  assign mesh_0_6_io_in_control_0_propagate = _T_392; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178936.4]
  assign mesh_0_6_io_in_control_0_shift = _T_390; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178926.4]
  assign mesh_0_6_io_in_valid_0 = _T_495_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179328.4]
  assign mesh_0_7_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177078.4]
  assign mesh_0_7_io_in_a_0 = _T_8_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177273.4]
  assign mesh_0_7_io_in_b_0 = {{11{_T_144_0[7]}},_T_144_0}; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177772.4]
  assign mesh_0_7_io_in_d_0 = {{11{_T_224_0[7]}},_T_224_0}; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@178124.4]
  assign mesh_0_7_io_in_control_0_propagate = _T_418; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@179062.4]
  assign mesh_0_7_io_in_control_0_shift = _T_416; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@179052.4]
  assign mesh_0_7_io_in_valid_0 = _T_504_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179354.4]
  assign mesh_1_0_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177081.4]
  assign mesh_1_0_io_in_a_0 = _T_10_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177278.4]
  assign mesh_1_0_io_in_b_0 = _T_75_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177469.4]
  assign mesh_1_0_io_in_d_0 = _T_155_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177821.4]
  assign mesh_1_0_io_in_control_0_propagate = _T_239; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178195.4]
  assign mesh_1_0_io_in_control_0_shift = _T_237; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178185.4]
  assign mesh_1_0_io_in_valid_0 = _T_442_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179175.4]
  assign mesh_1_1_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177084.4]
  assign mesh_1_1_io_in_a_0 = _T_11_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177281.4]
  assign mesh_1_1_io_in_b_0 = _T_85_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177513.4]
  assign mesh_1_1_io_in_d_0 = _T_165_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177865.4]
  assign mesh_1_1_io_in_control_0_propagate = _T_265; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178321.4]
  assign mesh_1_1_io_in_control_0_shift = _T_263; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178311.4]
  assign mesh_1_1_io_in_valid_0 = _T_451_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179201.4]
  assign mesh_1_2_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177087.4]
  assign mesh_1_2_io_in_a_0 = _T_12_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177284.4]
  assign mesh_1_2_io_in_b_0 = _T_95_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177557.4]
  assign mesh_1_2_io_in_d_0 = _T_175_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177909.4]
  assign mesh_1_2_io_in_control_0_propagate = _T_291; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178447.4]
  assign mesh_1_2_io_in_control_0_shift = _T_289; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178437.4]
  assign mesh_1_2_io_in_valid_0 = _T_460_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179227.4]
  assign mesh_1_3_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177090.4]
  assign mesh_1_3_io_in_a_0 = _T_13_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177287.4]
  assign mesh_1_3_io_in_b_0 = _T_105_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177601.4]
  assign mesh_1_3_io_in_d_0 = _T_185_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177953.4]
  assign mesh_1_3_io_in_control_0_propagate = _T_317; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178573.4]
  assign mesh_1_3_io_in_control_0_shift = _T_315; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178563.4]
  assign mesh_1_3_io_in_valid_0 = _T_469_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179253.4]
  assign mesh_1_4_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177093.4]
  assign mesh_1_4_io_in_a_0 = _T_14_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177290.4]
  assign mesh_1_4_io_in_b_0 = _T_115_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177645.4]
  assign mesh_1_4_io_in_d_0 = _T_195_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177997.4]
  assign mesh_1_4_io_in_control_0_propagate = _T_343; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178699.4]
  assign mesh_1_4_io_in_control_0_shift = _T_341; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178689.4]
  assign mesh_1_4_io_in_valid_0 = _T_478_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179279.4]
  assign mesh_1_5_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177096.4]
  assign mesh_1_5_io_in_a_0 = _T_15_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177293.4]
  assign mesh_1_5_io_in_b_0 = _T_125_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177689.4]
  assign mesh_1_5_io_in_d_0 = _T_205_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@178041.4]
  assign mesh_1_5_io_in_control_0_propagate = _T_369; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178825.4]
  assign mesh_1_5_io_in_control_0_shift = _T_367; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178815.4]
  assign mesh_1_5_io_in_valid_0 = _T_487_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179305.4]
  assign mesh_1_6_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177099.4]
  assign mesh_1_6_io_in_a_0 = _T_16_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177296.4]
  assign mesh_1_6_io_in_b_0 = _T_135_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177733.4]
  assign mesh_1_6_io_in_d_0 = _T_215_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@178085.4]
  assign mesh_1_6_io_in_control_0_propagate = _T_395; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178951.4]
  assign mesh_1_6_io_in_control_0_shift = _T_393; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178941.4]
  assign mesh_1_6_io_in_valid_0 = _T_496_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179331.4]
  assign mesh_1_7_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177102.4]
  assign mesh_1_7_io_in_a_0 = _T_17_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177299.4]
  assign mesh_1_7_io_in_b_0 = _T_145_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177777.4]
  assign mesh_1_7_io_in_d_0 = _T_225_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@178129.4]
  assign mesh_1_7_io_in_control_0_propagate = _T_421; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@179077.4]
  assign mesh_1_7_io_in_control_0_shift = _T_419; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@179067.4]
  assign mesh_1_7_io_in_valid_0 = _T_505_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179357.4]
  assign mesh_2_0_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177105.4]
  assign mesh_2_0_io_in_a_0 = _T_19_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177304.4]
  assign mesh_2_0_io_in_b_0 = _T_76_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177474.4]
  assign mesh_2_0_io_in_d_0 = _T_156_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177826.4]
  assign mesh_2_0_io_in_control_0_propagate = _T_242; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178210.4]
  assign mesh_2_0_io_in_control_0_shift = _T_240; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178200.4]
  assign mesh_2_0_io_in_valid_0 = _T_443_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179178.4]
  assign mesh_2_1_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177108.4]
  assign mesh_2_1_io_in_a_0 = _T_20_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177307.4]
  assign mesh_2_1_io_in_b_0 = _T_86_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177518.4]
  assign mesh_2_1_io_in_d_0 = _T_166_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177870.4]
  assign mesh_2_1_io_in_control_0_propagate = _T_268; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178336.4]
  assign mesh_2_1_io_in_control_0_shift = _T_266; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178326.4]
  assign mesh_2_1_io_in_valid_0 = _T_452_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179204.4]
  assign mesh_2_2_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177111.4]
  assign mesh_2_2_io_in_a_0 = _T_21_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177310.4]
  assign mesh_2_2_io_in_b_0 = _T_96_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177562.4]
  assign mesh_2_2_io_in_d_0 = _T_176_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177914.4]
  assign mesh_2_2_io_in_control_0_propagate = _T_294; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178462.4]
  assign mesh_2_2_io_in_control_0_shift = _T_292; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178452.4]
  assign mesh_2_2_io_in_valid_0 = _T_461_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179230.4]
  assign mesh_2_3_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177114.4]
  assign mesh_2_3_io_in_a_0 = _T_22_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177313.4]
  assign mesh_2_3_io_in_b_0 = _T_106_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177606.4]
  assign mesh_2_3_io_in_d_0 = _T_186_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177958.4]
  assign mesh_2_3_io_in_control_0_propagate = _T_320; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178588.4]
  assign mesh_2_3_io_in_control_0_shift = _T_318; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178578.4]
  assign mesh_2_3_io_in_valid_0 = _T_470_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179256.4]
  assign mesh_2_4_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177117.4]
  assign mesh_2_4_io_in_a_0 = _T_23_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177316.4]
  assign mesh_2_4_io_in_b_0 = _T_116_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177650.4]
  assign mesh_2_4_io_in_d_0 = _T_196_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@178002.4]
  assign mesh_2_4_io_in_control_0_propagate = _T_346; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178714.4]
  assign mesh_2_4_io_in_control_0_shift = _T_344; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178704.4]
  assign mesh_2_4_io_in_valid_0 = _T_479_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179282.4]
  assign mesh_2_5_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177120.4]
  assign mesh_2_5_io_in_a_0 = _T_24_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177319.4]
  assign mesh_2_5_io_in_b_0 = _T_126_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177694.4]
  assign mesh_2_5_io_in_d_0 = _T_206_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@178046.4]
  assign mesh_2_5_io_in_control_0_propagate = _T_372; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178840.4]
  assign mesh_2_5_io_in_control_0_shift = _T_370; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178830.4]
  assign mesh_2_5_io_in_valid_0 = _T_488_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179308.4]
  assign mesh_2_6_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177123.4]
  assign mesh_2_6_io_in_a_0 = _T_25_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177322.4]
  assign mesh_2_6_io_in_b_0 = _T_136_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177738.4]
  assign mesh_2_6_io_in_d_0 = _T_216_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@178090.4]
  assign mesh_2_6_io_in_control_0_propagate = _T_398; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178966.4]
  assign mesh_2_6_io_in_control_0_shift = _T_396; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178956.4]
  assign mesh_2_6_io_in_valid_0 = _T_497_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179334.4]
  assign mesh_2_7_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177126.4]
  assign mesh_2_7_io_in_a_0 = _T_26_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177325.4]
  assign mesh_2_7_io_in_b_0 = _T_146_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177782.4]
  assign mesh_2_7_io_in_d_0 = _T_226_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@178134.4]
  assign mesh_2_7_io_in_control_0_propagate = _T_424; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@179092.4]
  assign mesh_2_7_io_in_control_0_shift = _T_422; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@179082.4]
  assign mesh_2_7_io_in_valid_0 = _T_506_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179360.4]
  assign mesh_3_0_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177129.4]
  assign mesh_3_0_io_in_a_0 = _T_28_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177330.4]
  assign mesh_3_0_io_in_b_0 = _T_77_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177479.4]
  assign mesh_3_0_io_in_d_0 = _T_157_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177831.4]
  assign mesh_3_0_io_in_control_0_propagate = _T_245; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178225.4]
  assign mesh_3_0_io_in_control_0_shift = _T_243; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178215.4]
  assign mesh_3_0_io_in_valid_0 = _T_444_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179181.4]
  assign mesh_3_1_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177132.4]
  assign mesh_3_1_io_in_a_0 = _T_29_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177333.4]
  assign mesh_3_1_io_in_b_0 = _T_87_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177523.4]
  assign mesh_3_1_io_in_d_0 = _T_167_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177875.4]
  assign mesh_3_1_io_in_control_0_propagate = _T_271; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178351.4]
  assign mesh_3_1_io_in_control_0_shift = _T_269; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178341.4]
  assign mesh_3_1_io_in_valid_0 = _T_453_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179207.4]
  assign mesh_3_2_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177135.4]
  assign mesh_3_2_io_in_a_0 = _T_30_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177336.4]
  assign mesh_3_2_io_in_b_0 = _T_97_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177567.4]
  assign mesh_3_2_io_in_d_0 = _T_177_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177919.4]
  assign mesh_3_2_io_in_control_0_propagate = _T_297; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178477.4]
  assign mesh_3_2_io_in_control_0_shift = _T_295; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178467.4]
  assign mesh_3_2_io_in_valid_0 = _T_462_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179233.4]
  assign mesh_3_3_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177138.4]
  assign mesh_3_3_io_in_a_0 = _T_31_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177339.4]
  assign mesh_3_3_io_in_b_0 = _T_107_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177611.4]
  assign mesh_3_3_io_in_d_0 = _T_187_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177963.4]
  assign mesh_3_3_io_in_control_0_propagate = _T_323; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178603.4]
  assign mesh_3_3_io_in_control_0_shift = _T_321; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178593.4]
  assign mesh_3_3_io_in_valid_0 = _T_471_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179259.4]
  assign mesh_3_4_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177141.4]
  assign mesh_3_4_io_in_a_0 = _T_32_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177342.4]
  assign mesh_3_4_io_in_b_0 = _T_117_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177655.4]
  assign mesh_3_4_io_in_d_0 = _T_197_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@178007.4]
  assign mesh_3_4_io_in_control_0_propagate = _T_349; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178729.4]
  assign mesh_3_4_io_in_control_0_shift = _T_347; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178719.4]
  assign mesh_3_4_io_in_valid_0 = _T_480_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179285.4]
  assign mesh_3_5_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177144.4]
  assign mesh_3_5_io_in_a_0 = _T_33_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177345.4]
  assign mesh_3_5_io_in_b_0 = _T_127_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177699.4]
  assign mesh_3_5_io_in_d_0 = _T_207_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@178051.4]
  assign mesh_3_5_io_in_control_0_propagate = _T_375; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178855.4]
  assign mesh_3_5_io_in_control_0_shift = _T_373; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178845.4]
  assign mesh_3_5_io_in_valid_0 = _T_489_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179311.4]
  assign mesh_3_6_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177147.4]
  assign mesh_3_6_io_in_a_0 = _T_34_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177348.4]
  assign mesh_3_6_io_in_b_0 = _T_137_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177743.4]
  assign mesh_3_6_io_in_d_0 = _T_217_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@178095.4]
  assign mesh_3_6_io_in_control_0_propagate = _T_401; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178981.4]
  assign mesh_3_6_io_in_control_0_shift = _T_399; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178971.4]
  assign mesh_3_6_io_in_valid_0 = _T_498_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179337.4]
  assign mesh_3_7_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177150.4]
  assign mesh_3_7_io_in_a_0 = _T_35_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177351.4]
  assign mesh_3_7_io_in_b_0 = _T_147_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177787.4]
  assign mesh_3_7_io_in_d_0 = _T_227_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@178139.4]
  assign mesh_3_7_io_in_control_0_propagate = _T_427; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@179107.4]
  assign mesh_3_7_io_in_control_0_shift = _T_425; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@179097.4]
  assign mesh_3_7_io_in_valid_0 = _T_507_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179363.4]
  assign mesh_4_0_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177153.4]
  assign mesh_4_0_io_in_a_0 = _T_37_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177356.4]
  assign mesh_4_0_io_in_b_0 = _T_78_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177484.4]
  assign mesh_4_0_io_in_d_0 = _T_158_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177836.4]
  assign mesh_4_0_io_in_control_0_propagate = _T_248; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178240.4]
  assign mesh_4_0_io_in_control_0_shift = _T_246; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178230.4]
  assign mesh_4_0_io_in_valid_0 = _T_445_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179184.4]
  assign mesh_4_1_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177156.4]
  assign mesh_4_1_io_in_a_0 = _T_38_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177359.4]
  assign mesh_4_1_io_in_b_0 = _T_88_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177528.4]
  assign mesh_4_1_io_in_d_0 = _T_168_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177880.4]
  assign mesh_4_1_io_in_control_0_propagate = _T_274; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178366.4]
  assign mesh_4_1_io_in_control_0_shift = _T_272; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178356.4]
  assign mesh_4_1_io_in_valid_0 = _T_454_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179210.4]
  assign mesh_4_2_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177159.4]
  assign mesh_4_2_io_in_a_0 = _T_39_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177362.4]
  assign mesh_4_2_io_in_b_0 = _T_98_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177572.4]
  assign mesh_4_2_io_in_d_0 = _T_178_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177924.4]
  assign mesh_4_2_io_in_control_0_propagate = _T_300; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178492.4]
  assign mesh_4_2_io_in_control_0_shift = _T_298; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178482.4]
  assign mesh_4_2_io_in_valid_0 = _T_463_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179236.4]
  assign mesh_4_3_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177162.4]
  assign mesh_4_3_io_in_a_0 = _T_40_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177365.4]
  assign mesh_4_3_io_in_b_0 = _T_108_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177616.4]
  assign mesh_4_3_io_in_d_0 = _T_188_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177968.4]
  assign mesh_4_3_io_in_control_0_propagate = _T_326; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178618.4]
  assign mesh_4_3_io_in_control_0_shift = _T_324; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178608.4]
  assign mesh_4_3_io_in_valid_0 = _T_472_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179262.4]
  assign mesh_4_4_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177165.4]
  assign mesh_4_4_io_in_a_0 = _T_41_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177368.4]
  assign mesh_4_4_io_in_b_0 = _T_118_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177660.4]
  assign mesh_4_4_io_in_d_0 = _T_198_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@178012.4]
  assign mesh_4_4_io_in_control_0_propagate = _T_352; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178744.4]
  assign mesh_4_4_io_in_control_0_shift = _T_350; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178734.4]
  assign mesh_4_4_io_in_valid_0 = _T_481_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179288.4]
  assign mesh_4_5_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177168.4]
  assign mesh_4_5_io_in_a_0 = _T_42_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177371.4]
  assign mesh_4_5_io_in_b_0 = _T_128_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177704.4]
  assign mesh_4_5_io_in_d_0 = _T_208_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@178056.4]
  assign mesh_4_5_io_in_control_0_propagate = _T_378; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178870.4]
  assign mesh_4_5_io_in_control_0_shift = _T_376; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178860.4]
  assign mesh_4_5_io_in_valid_0 = _T_490_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179314.4]
  assign mesh_4_6_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177171.4]
  assign mesh_4_6_io_in_a_0 = _T_43_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177374.4]
  assign mesh_4_6_io_in_b_0 = _T_138_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177748.4]
  assign mesh_4_6_io_in_d_0 = _T_218_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@178100.4]
  assign mesh_4_6_io_in_control_0_propagate = _T_404; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178996.4]
  assign mesh_4_6_io_in_control_0_shift = _T_402; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178986.4]
  assign mesh_4_6_io_in_valid_0 = _T_499_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179340.4]
  assign mesh_4_7_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177174.4]
  assign mesh_4_7_io_in_a_0 = _T_44_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177377.4]
  assign mesh_4_7_io_in_b_0 = _T_148_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177792.4]
  assign mesh_4_7_io_in_d_0 = _T_228_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@178144.4]
  assign mesh_4_7_io_in_control_0_propagate = _T_430; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@179122.4]
  assign mesh_4_7_io_in_control_0_shift = _T_428; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@179112.4]
  assign mesh_4_7_io_in_valid_0 = _T_508_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179366.4]
  assign mesh_5_0_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177177.4]
  assign mesh_5_0_io_in_a_0 = _T_46_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177382.4]
  assign mesh_5_0_io_in_b_0 = _T_79_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177489.4]
  assign mesh_5_0_io_in_d_0 = _T_159_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177841.4]
  assign mesh_5_0_io_in_control_0_propagate = _T_251; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178255.4]
  assign mesh_5_0_io_in_control_0_shift = _T_249; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178245.4]
  assign mesh_5_0_io_in_valid_0 = _T_446_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179187.4]
  assign mesh_5_1_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177180.4]
  assign mesh_5_1_io_in_a_0 = _T_47_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177385.4]
  assign mesh_5_1_io_in_b_0 = _T_89_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177533.4]
  assign mesh_5_1_io_in_d_0 = _T_169_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177885.4]
  assign mesh_5_1_io_in_control_0_propagate = _T_277; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178381.4]
  assign mesh_5_1_io_in_control_0_shift = _T_275; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178371.4]
  assign mesh_5_1_io_in_valid_0 = _T_455_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179213.4]
  assign mesh_5_2_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177183.4]
  assign mesh_5_2_io_in_a_0 = _T_48_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177388.4]
  assign mesh_5_2_io_in_b_0 = _T_99_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177577.4]
  assign mesh_5_2_io_in_d_0 = _T_179_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177929.4]
  assign mesh_5_2_io_in_control_0_propagate = _T_303; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178507.4]
  assign mesh_5_2_io_in_control_0_shift = _T_301; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178497.4]
  assign mesh_5_2_io_in_valid_0 = _T_464_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179239.4]
  assign mesh_5_3_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177186.4]
  assign mesh_5_3_io_in_a_0 = _T_49_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177391.4]
  assign mesh_5_3_io_in_b_0 = _T_109_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177621.4]
  assign mesh_5_3_io_in_d_0 = _T_189_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177973.4]
  assign mesh_5_3_io_in_control_0_propagate = _T_329; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178633.4]
  assign mesh_5_3_io_in_control_0_shift = _T_327; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178623.4]
  assign mesh_5_3_io_in_valid_0 = _T_473_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179265.4]
  assign mesh_5_4_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177189.4]
  assign mesh_5_4_io_in_a_0 = _T_50_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177394.4]
  assign mesh_5_4_io_in_b_0 = _T_119_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177665.4]
  assign mesh_5_4_io_in_d_0 = _T_199_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@178017.4]
  assign mesh_5_4_io_in_control_0_propagate = _T_355; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178759.4]
  assign mesh_5_4_io_in_control_0_shift = _T_353; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178749.4]
  assign mesh_5_4_io_in_valid_0 = _T_482_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179291.4]
  assign mesh_5_5_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177192.4]
  assign mesh_5_5_io_in_a_0 = _T_51_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177397.4]
  assign mesh_5_5_io_in_b_0 = _T_129_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177709.4]
  assign mesh_5_5_io_in_d_0 = _T_209_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@178061.4]
  assign mesh_5_5_io_in_control_0_propagate = _T_381; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178885.4]
  assign mesh_5_5_io_in_control_0_shift = _T_379; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178875.4]
  assign mesh_5_5_io_in_valid_0 = _T_491_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179317.4]
  assign mesh_5_6_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177195.4]
  assign mesh_5_6_io_in_a_0 = _T_52_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177400.4]
  assign mesh_5_6_io_in_b_0 = _T_139_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177753.4]
  assign mesh_5_6_io_in_d_0 = _T_219_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@178105.4]
  assign mesh_5_6_io_in_control_0_propagate = _T_407; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@179011.4]
  assign mesh_5_6_io_in_control_0_shift = _T_405; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@179001.4]
  assign mesh_5_6_io_in_valid_0 = _T_500_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179343.4]
  assign mesh_5_7_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177198.4]
  assign mesh_5_7_io_in_a_0 = _T_53_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177403.4]
  assign mesh_5_7_io_in_b_0 = _T_149_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177797.4]
  assign mesh_5_7_io_in_d_0 = _T_229_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@178149.4]
  assign mesh_5_7_io_in_control_0_propagate = _T_433; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@179137.4]
  assign mesh_5_7_io_in_control_0_shift = _T_431; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@179127.4]
  assign mesh_5_7_io_in_valid_0 = _T_509_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179369.4]
  assign mesh_6_0_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177201.4]
  assign mesh_6_0_io_in_a_0 = _T_55_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177408.4]
  assign mesh_6_0_io_in_b_0 = _T_80_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177494.4]
  assign mesh_6_0_io_in_d_0 = _T_160_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177846.4]
  assign mesh_6_0_io_in_control_0_propagate = _T_254; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178270.4]
  assign mesh_6_0_io_in_control_0_shift = _T_252; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178260.4]
  assign mesh_6_0_io_in_valid_0 = _T_447_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179190.4]
  assign mesh_6_1_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177204.4]
  assign mesh_6_1_io_in_a_0 = _T_56_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177411.4]
  assign mesh_6_1_io_in_b_0 = _T_90_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177538.4]
  assign mesh_6_1_io_in_d_0 = _T_170_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177890.4]
  assign mesh_6_1_io_in_control_0_propagate = _T_280; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178396.4]
  assign mesh_6_1_io_in_control_0_shift = _T_278; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178386.4]
  assign mesh_6_1_io_in_valid_0 = _T_456_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179216.4]
  assign mesh_6_2_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177207.4]
  assign mesh_6_2_io_in_a_0 = _T_57_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177414.4]
  assign mesh_6_2_io_in_b_0 = _T_100_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177582.4]
  assign mesh_6_2_io_in_d_0 = _T_180_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177934.4]
  assign mesh_6_2_io_in_control_0_propagate = _T_306; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178522.4]
  assign mesh_6_2_io_in_control_0_shift = _T_304; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178512.4]
  assign mesh_6_2_io_in_valid_0 = _T_465_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179242.4]
  assign mesh_6_3_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177210.4]
  assign mesh_6_3_io_in_a_0 = _T_58_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177417.4]
  assign mesh_6_3_io_in_b_0 = _T_110_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177626.4]
  assign mesh_6_3_io_in_d_0 = _T_190_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177978.4]
  assign mesh_6_3_io_in_control_0_propagate = _T_332; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178648.4]
  assign mesh_6_3_io_in_control_0_shift = _T_330; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178638.4]
  assign mesh_6_3_io_in_valid_0 = _T_474_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179268.4]
  assign mesh_6_4_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177213.4]
  assign mesh_6_4_io_in_a_0 = _T_59_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177420.4]
  assign mesh_6_4_io_in_b_0 = _T_120_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177670.4]
  assign mesh_6_4_io_in_d_0 = _T_200_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@178022.4]
  assign mesh_6_4_io_in_control_0_propagate = _T_358; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178774.4]
  assign mesh_6_4_io_in_control_0_shift = _T_356; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178764.4]
  assign mesh_6_4_io_in_valid_0 = _T_483_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179294.4]
  assign mesh_6_5_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177216.4]
  assign mesh_6_5_io_in_a_0 = _T_60_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177423.4]
  assign mesh_6_5_io_in_b_0 = _T_130_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177714.4]
  assign mesh_6_5_io_in_d_0 = _T_210_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@178066.4]
  assign mesh_6_5_io_in_control_0_propagate = _T_384; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178900.4]
  assign mesh_6_5_io_in_control_0_shift = _T_382; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178890.4]
  assign mesh_6_5_io_in_valid_0 = _T_492_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179320.4]
  assign mesh_6_6_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177219.4]
  assign mesh_6_6_io_in_a_0 = _T_61_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177426.4]
  assign mesh_6_6_io_in_b_0 = _T_140_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177758.4]
  assign mesh_6_6_io_in_d_0 = _T_220_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@178110.4]
  assign mesh_6_6_io_in_control_0_propagate = _T_410; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@179026.4]
  assign mesh_6_6_io_in_control_0_shift = _T_408; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@179016.4]
  assign mesh_6_6_io_in_valid_0 = _T_501_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179346.4]
  assign mesh_6_7_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177222.4]
  assign mesh_6_7_io_in_a_0 = _T_62_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177429.4]
  assign mesh_6_7_io_in_b_0 = _T_150_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177802.4]
  assign mesh_6_7_io_in_d_0 = _T_230_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@178154.4]
  assign mesh_6_7_io_in_control_0_propagate = _T_436; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@179152.4]
  assign mesh_6_7_io_in_control_0_shift = _T_434; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@179142.4]
  assign mesh_6_7_io_in_valid_0 = _T_510_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179372.4]
  assign mesh_7_0_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177225.4]
  assign mesh_7_0_io_in_a_0 = _T_64_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177434.4]
  assign mesh_7_0_io_in_b_0 = _T_81_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177499.4]
  assign mesh_7_0_io_in_d_0 = _T_161_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177851.4]
  assign mesh_7_0_io_in_control_0_propagate = _T_257; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178285.4]
  assign mesh_7_0_io_in_control_0_shift = _T_255; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178275.4]
  assign mesh_7_0_io_in_valid_0 = _T_448_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179193.4]
  assign mesh_7_1_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177228.4]
  assign mesh_7_1_io_in_a_0 = _T_65_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177437.4]
  assign mesh_7_1_io_in_b_0 = _T_91_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177543.4]
  assign mesh_7_1_io_in_d_0 = _T_171_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177895.4]
  assign mesh_7_1_io_in_control_0_propagate = _T_283; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178411.4]
  assign mesh_7_1_io_in_control_0_shift = _T_281; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178401.4]
  assign mesh_7_1_io_in_valid_0 = _T_457_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179219.4]
  assign mesh_7_2_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177231.4]
  assign mesh_7_2_io_in_a_0 = _T_66_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177440.4]
  assign mesh_7_2_io_in_b_0 = _T_101_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177587.4]
  assign mesh_7_2_io_in_d_0 = _T_181_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177939.4]
  assign mesh_7_2_io_in_control_0_propagate = _T_309; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178537.4]
  assign mesh_7_2_io_in_control_0_shift = _T_307; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178527.4]
  assign mesh_7_2_io_in_valid_0 = _T_466_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179245.4]
  assign mesh_7_3_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177234.4]
  assign mesh_7_3_io_in_a_0 = _T_67_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177443.4]
  assign mesh_7_3_io_in_b_0 = _T_111_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177631.4]
  assign mesh_7_3_io_in_d_0 = _T_191_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177983.4]
  assign mesh_7_3_io_in_control_0_propagate = _T_335; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178663.4]
  assign mesh_7_3_io_in_control_0_shift = _T_333; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178653.4]
  assign mesh_7_3_io_in_valid_0 = _T_475_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179271.4]
  assign mesh_7_4_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177237.4]
  assign mesh_7_4_io_in_a_0 = _T_68_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177446.4]
  assign mesh_7_4_io_in_b_0 = _T_121_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177675.4]
  assign mesh_7_4_io_in_d_0 = _T_201_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@178027.4]
  assign mesh_7_4_io_in_control_0_propagate = _T_361; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178789.4]
  assign mesh_7_4_io_in_control_0_shift = _T_359; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178779.4]
  assign mesh_7_4_io_in_valid_0 = _T_484_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179297.4]
  assign mesh_7_5_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177240.4]
  assign mesh_7_5_io_in_a_0 = _T_69_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177449.4]
  assign mesh_7_5_io_in_b_0 = _T_131_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177719.4]
  assign mesh_7_5_io_in_d_0 = _T_211_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@178071.4]
  assign mesh_7_5_io_in_control_0_propagate = _T_387; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@178915.4]
  assign mesh_7_5_io_in_control_0_shift = _T_385; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@178905.4]
  assign mesh_7_5_io_in_valid_0 = _T_493_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179323.4]
  assign mesh_7_6_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177243.4]
  assign mesh_7_6_io_in_a_0 = _T_70_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177452.4]
  assign mesh_7_6_io_in_b_0 = _T_141_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177763.4]
  assign mesh_7_6_io_in_d_0 = _T_221_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@178115.4]
  assign mesh_7_6_io_in_control_0_propagate = _T_413; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@179041.4]
  assign mesh_7_6_io_in_control_0_shift = _T_411; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@179031.4]
  assign mesh_7_6_io_in_valid_0 = _T_502_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179349.4]
  assign mesh_7_7_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig.fir@177246.4]
  assign mesh_7_7_io_in_a_0 = _T_71_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177455.4]
  assign mesh_7_7_io_in_b_0 = _T_151_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@177807.4]
  assign mesh_7_7_io_in_d_0 = _T_231_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig.fir@178159.4]
  assign mesh_7_7_io_in_control_0_propagate = _T_439; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig.fir@179167.4]
  assign mesh_7_7_io_in_control_0_shift = _T_437; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig.fir@179157.4]
  assign mesh_7_7_io_in_valid_0 = _T_511_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig.fir@179375.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_0 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1_0 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2_0 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_3_0 = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_4_0 = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_5_0 = _RAND_5[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_6_0 = _RAND_6[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_7_0 = _RAND_7[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_8_0 = _RAND_8[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_9_0 = _RAND_9[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_10_0 = _RAND_10[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_11_0 = _RAND_11[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_12_0 = _RAND_12[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_13_0 = _RAND_13[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_14_0 = _RAND_14[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_15_0 = _RAND_15[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_16_0 = _RAND_16[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_17_0 = _RAND_17[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_18_0 = _RAND_18[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_19_0 = _RAND_19[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_20_0 = _RAND_20[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_21_0 = _RAND_21[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_22_0 = _RAND_22[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_23_0 = _RAND_23[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_24_0 = _RAND_24[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_25_0 = _RAND_25[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_26_0 = _RAND_26[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_27_0 = _RAND_27[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_28_0 = _RAND_28[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_29_0 = _RAND_29[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_30_0 = _RAND_30[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_31_0 = _RAND_31[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_32_0 = _RAND_32[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_33_0 = _RAND_33[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_34_0 = _RAND_34[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_35_0 = _RAND_35[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_36_0 = _RAND_36[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_37_0 = _RAND_37[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_38_0 = _RAND_38[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_39_0 = _RAND_39[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_40_0 = _RAND_40[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_41_0 = _RAND_41[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_42_0 = _RAND_42[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_43_0 = _RAND_43[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_44_0 = _RAND_44[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_45_0 = _RAND_45[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_46_0 = _RAND_46[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_47_0 = _RAND_47[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_48_0 = _RAND_48[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_49_0 = _RAND_49[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_50_0 = _RAND_50[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_51_0 = _RAND_51[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_52_0 = _RAND_52[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_53_0 = _RAND_53[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_54_0 = _RAND_54[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_55_0 = _RAND_55[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_56_0 = _RAND_56[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_57_0 = _RAND_57[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_58_0 = _RAND_58[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_59_0 = _RAND_59[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_60_0 = _RAND_60[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_61_0 = _RAND_61[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_62_0 = _RAND_62[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_63_0 = _RAND_63[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_64_0 = _RAND_64[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_65_0 = _RAND_65[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_66_0 = _RAND_66[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_67_0 = _RAND_67[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_68_0 = _RAND_68[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_69_0 = _RAND_69[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_70_0 = _RAND_70[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_71_0 = _RAND_71[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_72_0 = _RAND_72[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_73_0 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_74_0 = _RAND_74[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_75_0 = _RAND_75[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_76_0 = _RAND_76[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_77_0 = _RAND_77[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_78_0 = _RAND_78[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_79_0 = _RAND_79[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_80_0 = _RAND_80[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_81_0 = _RAND_81[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_82_0 = _RAND_82[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_83_0 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_84_0 = _RAND_84[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_85_0 = _RAND_85[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_86_0 = _RAND_86[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_87_0 = _RAND_87[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_88_0 = _RAND_88[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_89_0 = _RAND_89[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_90_0 = _RAND_90[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_91_0 = _RAND_91[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_92_0 = _RAND_92[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_93_0 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_94_0 = _RAND_94[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_95_0 = _RAND_95[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_96_0 = _RAND_96[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_97_0 = _RAND_97[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_98_0 = _RAND_98[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_99_0 = _RAND_99[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_100_0 = _RAND_100[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_101_0 = _RAND_101[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_102_0 = _RAND_102[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_103_0 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_104_0 = _RAND_104[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_105_0 = _RAND_105[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_106_0 = _RAND_106[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_107_0 = _RAND_107[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_108_0 = _RAND_108[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_109_0 = _RAND_109[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_110_0 = _RAND_110[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_111_0 = _RAND_111[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_112_0 = _RAND_112[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_113_0 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_114_0 = _RAND_114[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_115_0 = _RAND_115[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_116_0 = _RAND_116[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_117_0 = _RAND_117[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_118_0 = _RAND_118[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_119_0 = _RAND_119[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_120_0 = _RAND_120[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_121_0 = _RAND_121[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_122_0 = _RAND_122[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_123_0 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_124_0 = _RAND_124[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_125_0 = _RAND_125[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_126_0 = _RAND_126[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_127_0 = _RAND_127[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_128_0 = _RAND_128[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_129_0 = _RAND_129[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T_130_0 = _RAND_130[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _T_131_0 = _RAND_131[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _T_132_0 = _RAND_132[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _T_133_0 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T_134_0 = _RAND_134[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _T_135_0 = _RAND_135[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _T_136_0 = _RAND_136[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _T_137_0 = _RAND_137[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T_138_0 = _RAND_138[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T_139_0 = _RAND_139[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _T_140_0 = _RAND_140[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _T_141_0 = _RAND_141[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T_142_0 = _RAND_142[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T_143_0 = _RAND_143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _T_144_0 = _RAND_144[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T_145_0 = _RAND_145[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T_146_0 = _RAND_146[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _T_147_0 = _RAND_147[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _T_148_0 = _RAND_148[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _T_149_0 = _RAND_149[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _T_150_0 = _RAND_150[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _T_151_0 = _RAND_151[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _T_152_0 = _RAND_152[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _T_153_0 = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T_154_0 = _RAND_154[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T_155_0 = _RAND_155[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T_156_0 = _RAND_156[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T_157_0 = _RAND_157[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T_158_0 = _RAND_158[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _T_159_0 = _RAND_159[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _T_160_0 = _RAND_160[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _T_161_0 = _RAND_161[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T_162_0 = _RAND_162[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T_163_0 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _T_164_0 = _RAND_164[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _T_165_0 = _RAND_165[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _T_166_0 = _RAND_166[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _T_167_0 = _RAND_167[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _T_168_0 = _RAND_168[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _T_169_0 = _RAND_169[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _T_170_0 = _RAND_170[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _T_171_0 = _RAND_171[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _T_172_0 = _RAND_172[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _T_173_0 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _T_174_0 = _RAND_174[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _T_175_0 = _RAND_175[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _T_176_0 = _RAND_176[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _T_177_0 = _RAND_177[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _T_178_0 = _RAND_178[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _T_179_0 = _RAND_179[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _T_180_0 = _RAND_180[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _T_181_0 = _RAND_181[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _T_182_0 = _RAND_182[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _T_183_0 = _RAND_183[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T_184_0 = _RAND_184[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _T_185_0 = _RAND_185[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _T_186_0 = _RAND_186[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _T_187_0 = _RAND_187[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _T_188_0 = _RAND_188[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _T_189_0 = _RAND_189[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T_190_0 = _RAND_190[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _T_191_0 = _RAND_191[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _T_192_0 = _RAND_192[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _T_193_0 = _RAND_193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _T_194_0 = _RAND_194[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _T_195_0 = _RAND_195[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _T_196_0 = _RAND_196[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _T_197_0 = _RAND_197[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _T_198_0 = _RAND_198[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _T_199_0 = _RAND_199[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _T_200_0 = _RAND_200[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _T_201_0 = _RAND_201[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _T_202_0 = _RAND_202[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _T_203_0 = _RAND_203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _T_204_0 = _RAND_204[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _T_205_0 = _RAND_205[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _T_206_0 = _RAND_206[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _T_207_0 = _RAND_207[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _T_208_0 = _RAND_208[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _T_209_0 = _RAND_209[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _T_210_0 = _RAND_210[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _T_211_0 = _RAND_211[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _T_212_0 = _RAND_212[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _T_213_0 = _RAND_213[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _T_214_0 = _RAND_214[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _T_215_0 = _RAND_215[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _T_216_0 = _RAND_216[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _T_217_0 = _RAND_217[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _T_218_0 = _RAND_218[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _T_219_0 = _RAND_219[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _T_220_0 = _RAND_220[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _T_221_0 = _RAND_221[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _T_222_0 = _RAND_222[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _T_223_0 = _RAND_223[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  _T_224_0 = _RAND_224[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  _T_225_0 = _RAND_225[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  _T_226_0 = _RAND_226[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  _T_227_0 = _RAND_227[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  _T_228_0 = _RAND_228[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  _T_229_0 = _RAND_229[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  _T_230_0 = _RAND_230[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  _T_231_0 = _RAND_231[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  _T_232_0_propagate = _RAND_232[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  _T_232_0_shift = _RAND_233[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  _T_233_0 = _RAND_234[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  _T_234 = _RAND_235[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  _T_236 = _RAND_236[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  _T_237 = _RAND_237[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  _T_239 = _RAND_238[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  _T_240 = _RAND_239[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  _T_242 = _RAND_240[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  _T_243 = _RAND_241[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  _T_245 = _RAND_242[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  _T_246 = _RAND_243[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  _T_248 = _RAND_244[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  _T_249 = _RAND_245[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  _T_251 = _RAND_246[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  _T_252 = _RAND_247[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  _T_254 = _RAND_248[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  _T_255 = _RAND_249[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  _T_257 = _RAND_250[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  _T_258_0_propagate = _RAND_251[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  _T_258_0_shift = _RAND_252[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  _T_259_0 = _RAND_253[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _T_260 = _RAND_254[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _T_262 = _RAND_255[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  _T_263 = _RAND_256[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  _T_265 = _RAND_257[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  _T_266 = _RAND_258[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  _T_268 = _RAND_259[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  _T_269 = _RAND_260[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  _T_271 = _RAND_261[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  _T_272 = _RAND_262[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  _T_274 = _RAND_263[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  _T_275 = _RAND_264[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  _T_277 = _RAND_265[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  _T_278 = _RAND_266[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  _T_280 = _RAND_267[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  _T_281 = _RAND_268[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  _T_283 = _RAND_269[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  _T_284_0_propagate = _RAND_270[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  _T_284_0_shift = _RAND_271[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  _T_285_0 = _RAND_272[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  _T_286 = _RAND_273[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  _T_288 = _RAND_274[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  _T_289 = _RAND_275[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  _T_291 = _RAND_276[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  _T_292 = _RAND_277[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  _T_294 = _RAND_278[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  _T_295 = _RAND_279[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  _T_297 = _RAND_280[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  _T_298 = _RAND_281[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  _T_300 = _RAND_282[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  _T_301 = _RAND_283[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  _T_303 = _RAND_284[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  _T_304 = _RAND_285[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  _T_306 = _RAND_286[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  _T_307 = _RAND_287[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  _T_309 = _RAND_288[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  _T_310_0_propagate = _RAND_289[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  _T_310_0_shift = _RAND_290[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  _T_311_0 = _RAND_291[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  _T_312 = _RAND_292[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  _T_314 = _RAND_293[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  _T_315 = _RAND_294[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  _T_317 = _RAND_295[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  _T_318 = _RAND_296[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  _T_320 = _RAND_297[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  _T_321 = _RAND_298[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  _T_323 = _RAND_299[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  _T_324 = _RAND_300[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  _T_326 = _RAND_301[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  _T_327 = _RAND_302[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  _T_329 = _RAND_303[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  _T_330 = _RAND_304[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  _T_332 = _RAND_305[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  _T_333 = _RAND_306[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  _T_335 = _RAND_307[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  _T_336_0_propagate = _RAND_308[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  _T_336_0_shift = _RAND_309[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  _T_337_0 = _RAND_310[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  _T_338 = _RAND_311[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  _T_340 = _RAND_312[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  _T_341 = _RAND_313[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  _T_343 = _RAND_314[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  _T_344 = _RAND_315[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  _T_346 = _RAND_316[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  _T_347 = _RAND_317[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  _T_349 = _RAND_318[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  _T_350 = _RAND_319[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  _T_352 = _RAND_320[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  _T_353 = _RAND_321[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  _T_355 = _RAND_322[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  _T_356 = _RAND_323[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  _T_358 = _RAND_324[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  _T_359 = _RAND_325[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  _T_361 = _RAND_326[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  _T_362_0_propagate = _RAND_327[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  _T_362_0_shift = _RAND_328[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  _T_363_0 = _RAND_329[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  _T_364 = _RAND_330[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  _T_366 = _RAND_331[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  _T_367 = _RAND_332[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  _T_369 = _RAND_333[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  _T_370 = _RAND_334[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  _T_372 = _RAND_335[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  _T_373 = _RAND_336[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  _T_375 = _RAND_337[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  _T_376 = _RAND_338[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  _T_378 = _RAND_339[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  _T_379 = _RAND_340[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  _T_381 = _RAND_341[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  _T_382 = _RAND_342[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  _T_384 = _RAND_343[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  _T_385 = _RAND_344[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  _T_387 = _RAND_345[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  _T_388_0_propagate = _RAND_346[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  _T_388_0_shift = _RAND_347[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  _T_389_0 = _RAND_348[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  _T_390 = _RAND_349[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  _T_392 = _RAND_350[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  _T_393 = _RAND_351[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  _T_395 = _RAND_352[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  _T_396 = _RAND_353[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  _T_398 = _RAND_354[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  _T_399 = _RAND_355[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  _T_401 = _RAND_356[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  _T_402 = _RAND_357[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  _T_404 = _RAND_358[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  _T_405 = _RAND_359[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  _T_407 = _RAND_360[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  _T_408 = _RAND_361[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  _T_410 = _RAND_362[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  _T_411 = _RAND_363[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  _T_413 = _RAND_364[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  _T_414_0_propagate = _RAND_365[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  _T_414_0_shift = _RAND_366[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  _T_415_0 = _RAND_367[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  _T_416 = _RAND_368[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  _T_418 = _RAND_369[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  _T_419 = _RAND_370[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  _T_421 = _RAND_371[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  _T_422 = _RAND_372[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  _T_424 = _RAND_373[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  _T_425 = _RAND_374[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  _T_427 = _RAND_375[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  _T_428 = _RAND_376[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  _T_430 = _RAND_377[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  _T_431 = _RAND_378[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  _T_433 = _RAND_379[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  _T_434 = _RAND_380[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  _T_436 = _RAND_381[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  _T_437 = _RAND_382[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  _T_439 = _RAND_383[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  _T_440_0 = _RAND_384[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  _T_441_0 = _RAND_385[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  _T_442_0 = _RAND_386[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  _T_443_0 = _RAND_387[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  _T_444_0 = _RAND_388[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  _T_445_0 = _RAND_389[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  _T_446_0 = _RAND_390[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  _T_447_0 = _RAND_391[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  _T_448_0 = _RAND_392[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  _T_449_0 = _RAND_393[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  _T_450_0 = _RAND_394[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  _T_451_0 = _RAND_395[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  _T_452_0 = _RAND_396[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  _T_453_0 = _RAND_397[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  _T_454_0 = _RAND_398[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  _T_455_0 = _RAND_399[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{`RANDOM}};
  _T_456_0 = _RAND_400[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{`RANDOM}};
  _T_457_0 = _RAND_401[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{`RANDOM}};
  _T_458_0 = _RAND_402[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{`RANDOM}};
  _T_459_0 = _RAND_403[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{`RANDOM}};
  _T_460_0 = _RAND_404[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{`RANDOM}};
  _T_461_0 = _RAND_405[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{`RANDOM}};
  _T_462_0 = _RAND_406[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{`RANDOM}};
  _T_463_0 = _RAND_407[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {1{`RANDOM}};
  _T_464_0 = _RAND_408[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {1{`RANDOM}};
  _T_465_0 = _RAND_409[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {1{`RANDOM}};
  _T_466_0 = _RAND_410[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {1{`RANDOM}};
  _T_467_0 = _RAND_411[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {1{`RANDOM}};
  _T_468_0 = _RAND_412[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {1{`RANDOM}};
  _T_469_0 = _RAND_413[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {1{`RANDOM}};
  _T_470_0 = _RAND_414[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {1{`RANDOM}};
  _T_471_0 = _RAND_415[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {1{`RANDOM}};
  _T_472_0 = _RAND_416[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {1{`RANDOM}};
  _T_473_0 = _RAND_417[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {1{`RANDOM}};
  _T_474_0 = _RAND_418[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {1{`RANDOM}};
  _T_475_0 = _RAND_419[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {1{`RANDOM}};
  _T_476_0 = _RAND_420[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {1{`RANDOM}};
  _T_477_0 = _RAND_421[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {1{`RANDOM}};
  _T_478_0 = _RAND_422[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {1{`RANDOM}};
  _T_479_0 = _RAND_423[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {1{`RANDOM}};
  _T_480_0 = _RAND_424[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {1{`RANDOM}};
  _T_481_0 = _RAND_425[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {1{`RANDOM}};
  _T_482_0 = _RAND_426[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {1{`RANDOM}};
  _T_483_0 = _RAND_427[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {1{`RANDOM}};
  _T_484_0 = _RAND_428[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {1{`RANDOM}};
  _T_485_0 = _RAND_429[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {1{`RANDOM}};
  _T_486_0 = _RAND_430[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {1{`RANDOM}};
  _T_487_0 = _RAND_431[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {1{`RANDOM}};
  _T_488_0 = _RAND_432[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {1{`RANDOM}};
  _T_489_0 = _RAND_433[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {1{`RANDOM}};
  _T_490_0 = _RAND_434[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {1{`RANDOM}};
  _T_491_0 = _RAND_435[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {1{`RANDOM}};
  _T_492_0 = _RAND_436[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {1{`RANDOM}};
  _T_493_0 = _RAND_437[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {1{`RANDOM}};
  _T_494_0 = _RAND_438[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {1{`RANDOM}};
  _T_495_0 = _RAND_439[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {1{`RANDOM}};
  _T_496_0 = _RAND_440[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {1{`RANDOM}};
  _T_497_0 = _RAND_441[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {1{`RANDOM}};
  _T_498_0 = _RAND_442[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_443 = {1{`RANDOM}};
  _T_499_0 = _RAND_443[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_444 = {1{`RANDOM}};
  _T_500_0 = _RAND_444[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_445 = {1{`RANDOM}};
  _T_501_0 = _RAND_445[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_446 = {1{`RANDOM}};
  _T_502_0 = _RAND_446[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_447 = {1{`RANDOM}};
  _T_503_0 = _RAND_447[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_448 = {1{`RANDOM}};
  _T_504_0 = _RAND_448[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_449 = {1{`RANDOM}};
  _T_505_0 = _RAND_449[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_450 = {1{`RANDOM}};
  _T_506_0 = _RAND_450[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_451 = {1{`RANDOM}};
  _T_507_0 = _RAND_451[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_452 = {1{`RANDOM}};
  _T_508_0 = _RAND_452[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_453 = {1{`RANDOM}};
  _T_509_0 = _RAND_453[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_454 = {1{`RANDOM}};
  _T_510_0 = _RAND_454[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_455 = {1{`RANDOM}};
  _T_511_0 = _RAND_455[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    _T_0 <= io_in_a_0_0;
    _T_1_0 <= _T_0;
    _T_2_0 <= mesh_0_0_io_out_a_0;
    _T_3_0 <= mesh_0_1_io_out_a_0;
    _T_4_0 <= mesh_0_2_io_out_a_0;
    _T_5_0 <= mesh_0_3_io_out_a_0;
    _T_6_0 <= mesh_0_4_io_out_a_0;
    _T_7_0 <= mesh_0_5_io_out_a_0;
    _T_8_0 <= mesh_0_6_io_out_a_0;
    _T_9_0 <= io_in_a_1_0;
    _T_10_0 <= _T_9_0;
    _T_11_0 <= mesh_1_0_io_out_a_0;
    _T_12_0 <= mesh_1_1_io_out_a_0;
    _T_13_0 <= mesh_1_2_io_out_a_0;
    _T_14_0 <= mesh_1_3_io_out_a_0;
    _T_15_0 <= mesh_1_4_io_out_a_0;
    _T_16_0 <= mesh_1_5_io_out_a_0;
    _T_17_0 <= mesh_1_6_io_out_a_0;
    _T_18_0 <= io_in_a_2_0;
    _T_19_0 <= _T_18_0;
    _T_20_0 <= mesh_2_0_io_out_a_0;
    _T_21_0 <= mesh_2_1_io_out_a_0;
    _T_22_0 <= mesh_2_2_io_out_a_0;
    _T_23_0 <= mesh_2_3_io_out_a_0;
    _T_24_0 <= mesh_2_4_io_out_a_0;
    _T_25_0 <= mesh_2_5_io_out_a_0;
    _T_26_0 <= mesh_2_6_io_out_a_0;
    _T_27_0 <= io_in_a_3_0;
    _T_28_0 <= _T_27_0;
    _T_29_0 <= mesh_3_0_io_out_a_0;
    _T_30_0 <= mesh_3_1_io_out_a_0;
    _T_31_0 <= mesh_3_2_io_out_a_0;
    _T_32_0 <= mesh_3_3_io_out_a_0;
    _T_33_0 <= mesh_3_4_io_out_a_0;
    _T_34_0 <= mesh_3_5_io_out_a_0;
    _T_35_0 <= mesh_3_6_io_out_a_0;
    _T_36_0 <= io_in_a_4_0;
    _T_37_0 <= _T_36_0;
    _T_38_0 <= mesh_4_0_io_out_a_0;
    _T_39_0 <= mesh_4_1_io_out_a_0;
    _T_40_0 <= mesh_4_2_io_out_a_0;
    _T_41_0 <= mesh_4_3_io_out_a_0;
    _T_42_0 <= mesh_4_4_io_out_a_0;
    _T_43_0 <= mesh_4_5_io_out_a_0;
    _T_44_0 <= mesh_4_6_io_out_a_0;
    _T_45_0 <= io_in_a_5_0;
    _T_46_0 <= _T_45_0;
    _T_47_0 <= mesh_5_0_io_out_a_0;
    _T_48_0 <= mesh_5_1_io_out_a_0;
    _T_49_0 <= mesh_5_2_io_out_a_0;
    _T_50_0 <= mesh_5_3_io_out_a_0;
    _T_51_0 <= mesh_5_4_io_out_a_0;
    _T_52_0 <= mesh_5_5_io_out_a_0;
    _T_53_0 <= mesh_5_6_io_out_a_0;
    _T_54_0 <= io_in_a_6_0;
    _T_55_0 <= _T_54_0;
    _T_56_0 <= mesh_6_0_io_out_a_0;
    _T_57_0 <= mesh_6_1_io_out_a_0;
    _T_58_0 <= mesh_6_2_io_out_a_0;
    _T_59_0 <= mesh_6_3_io_out_a_0;
    _T_60_0 <= mesh_6_4_io_out_a_0;
    _T_61_0 <= mesh_6_5_io_out_a_0;
    _T_62_0 <= mesh_6_6_io_out_a_0;
    _T_63_0 <= io_in_a_7_0;
    _T_64_0 <= _T_63_0;
    _T_65_0 <= mesh_7_0_io_out_a_0;
    _T_66_0 <= mesh_7_1_io_out_a_0;
    _T_67_0 <= mesh_7_2_io_out_a_0;
    _T_68_0 <= mesh_7_3_io_out_a_0;
    _T_69_0 <= mesh_7_4_io_out_a_0;
    _T_70_0 <= mesh_7_5_io_out_a_0;
    _T_71_0 <= mesh_7_6_io_out_a_0;
    _T_72_0 <= io_in_d_0_0;
    _T_73_0 <= io_in_valid_0_0;
    if (_T_73_0) begin
      _T_74_0 <= _T_72_0;
    end
    if (mesh_0_0_io_out_valid_0) begin
      _T_75_0 <= mesh_0_0_io_out_b_0;
    end
    if (mesh_1_0_io_out_valid_0) begin
      _T_76_0 <= mesh_1_0_io_out_b_0;
    end
    if (mesh_2_0_io_out_valid_0) begin
      _T_77_0 <= mesh_2_0_io_out_b_0;
    end
    if (mesh_3_0_io_out_valid_0) begin
      _T_78_0 <= mesh_3_0_io_out_b_0;
    end
    if (mesh_4_0_io_out_valid_0) begin
      _T_79_0 <= mesh_4_0_io_out_b_0;
    end
    if (mesh_5_0_io_out_valid_0) begin
      _T_80_0 <= mesh_5_0_io_out_b_0;
    end
    if (mesh_6_0_io_out_valid_0) begin
      _T_81_0 <= mesh_6_0_io_out_b_0;
    end
    _T_82_0 <= io_in_d_1_0;
    _T_83_0 <= io_in_valid_1_0;
    if (_T_83_0) begin
      _T_84_0 <= _T_82_0;
    end
    if (mesh_0_1_io_out_valid_0) begin
      _T_85_0 <= mesh_0_1_io_out_b_0;
    end
    if (mesh_1_1_io_out_valid_0) begin
      _T_86_0 <= mesh_1_1_io_out_b_0;
    end
    if (mesh_2_1_io_out_valid_0) begin
      _T_87_0 <= mesh_2_1_io_out_b_0;
    end
    if (mesh_3_1_io_out_valid_0) begin
      _T_88_0 <= mesh_3_1_io_out_b_0;
    end
    if (mesh_4_1_io_out_valid_0) begin
      _T_89_0 <= mesh_4_1_io_out_b_0;
    end
    if (mesh_5_1_io_out_valid_0) begin
      _T_90_0 <= mesh_5_1_io_out_b_0;
    end
    if (mesh_6_1_io_out_valid_0) begin
      _T_91_0 <= mesh_6_1_io_out_b_0;
    end
    _T_92_0 <= io_in_d_2_0;
    _T_93_0 <= io_in_valid_2_0;
    if (_T_93_0) begin
      _T_94_0 <= _T_92_0;
    end
    if (mesh_0_2_io_out_valid_0) begin
      _T_95_0 <= mesh_0_2_io_out_b_0;
    end
    if (mesh_1_2_io_out_valid_0) begin
      _T_96_0 <= mesh_1_2_io_out_b_0;
    end
    if (mesh_2_2_io_out_valid_0) begin
      _T_97_0 <= mesh_2_2_io_out_b_0;
    end
    if (mesh_3_2_io_out_valid_0) begin
      _T_98_0 <= mesh_3_2_io_out_b_0;
    end
    if (mesh_4_2_io_out_valid_0) begin
      _T_99_0 <= mesh_4_2_io_out_b_0;
    end
    if (mesh_5_2_io_out_valid_0) begin
      _T_100_0 <= mesh_5_2_io_out_b_0;
    end
    if (mesh_6_2_io_out_valid_0) begin
      _T_101_0 <= mesh_6_2_io_out_b_0;
    end
    _T_102_0 <= io_in_d_3_0;
    _T_103_0 <= io_in_valid_3_0;
    if (_T_103_0) begin
      _T_104_0 <= _T_102_0;
    end
    if (mesh_0_3_io_out_valid_0) begin
      _T_105_0 <= mesh_0_3_io_out_b_0;
    end
    if (mesh_1_3_io_out_valid_0) begin
      _T_106_0 <= mesh_1_3_io_out_b_0;
    end
    if (mesh_2_3_io_out_valid_0) begin
      _T_107_0 <= mesh_2_3_io_out_b_0;
    end
    if (mesh_3_3_io_out_valid_0) begin
      _T_108_0 <= mesh_3_3_io_out_b_0;
    end
    if (mesh_4_3_io_out_valid_0) begin
      _T_109_0 <= mesh_4_3_io_out_b_0;
    end
    if (mesh_5_3_io_out_valid_0) begin
      _T_110_0 <= mesh_5_3_io_out_b_0;
    end
    if (mesh_6_3_io_out_valid_0) begin
      _T_111_0 <= mesh_6_3_io_out_b_0;
    end
    _T_112_0 <= io_in_d_4_0;
    _T_113_0 <= io_in_valid_4_0;
    if (_T_113_0) begin
      _T_114_0 <= _T_112_0;
    end
    if (mesh_0_4_io_out_valid_0) begin
      _T_115_0 <= mesh_0_4_io_out_b_0;
    end
    if (mesh_1_4_io_out_valid_0) begin
      _T_116_0 <= mesh_1_4_io_out_b_0;
    end
    if (mesh_2_4_io_out_valid_0) begin
      _T_117_0 <= mesh_2_4_io_out_b_0;
    end
    if (mesh_3_4_io_out_valid_0) begin
      _T_118_0 <= mesh_3_4_io_out_b_0;
    end
    if (mesh_4_4_io_out_valid_0) begin
      _T_119_0 <= mesh_4_4_io_out_b_0;
    end
    if (mesh_5_4_io_out_valid_0) begin
      _T_120_0 <= mesh_5_4_io_out_b_0;
    end
    if (mesh_6_4_io_out_valid_0) begin
      _T_121_0 <= mesh_6_4_io_out_b_0;
    end
    _T_122_0 <= io_in_d_5_0;
    _T_123_0 <= io_in_valid_5_0;
    if (_T_123_0) begin
      _T_124_0 <= _T_122_0;
    end
    if (mesh_0_5_io_out_valid_0) begin
      _T_125_0 <= mesh_0_5_io_out_b_0;
    end
    if (mesh_1_5_io_out_valid_0) begin
      _T_126_0 <= mesh_1_5_io_out_b_0;
    end
    if (mesh_2_5_io_out_valid_0) begin
      _T_127_0 <= mesh_2_5_io_out_b_0;
    end
    if (mesh_3_5_io_out_valid_0) begin
      _T_128_0 <= mesh_3_5_io_out_b_0;
    end
    if (mesh_4_5_io_out_valid_0) begin
      _T_129_0 <= mesh_4_5_io_out_b_0;
    end
    if (mesh_5_5_io_out_valid_0) begin
      _T_130_0 <= mesh_5_5_io_out_b_0;
    end
    if (mesh_6_5_io_out_valid_0) begin
      _T_131_0 <= mesh_6_5_io_out_b_0;
    end
    _T_132_0 <= io_in_d_6_0;
    _T_133_0 <= io_in_valid_6_0;
    if (_T_133_0) begin
      _T_134_0 <= _T_132_0;
    end
    if (mesh_0_6_io_out_valid_0) begin
      _T_135_0 <= mesh_0_6_io_out_b_0;
    end
    if (mesh_1_6_io_out_valid_0) begin
      _T_136_0 <= mesh_1_6_io_out_b_0;
    end
    if (mesh_2_6_io_out_valid_0) begin
      _T_137_0 <= mesh_2_6_io_out_b_0;
    end
    if (mesh_3_6_io_out_valid_0) begin
      _T_138_0 <= mesh_3_6_io_out_b_0;
    end
    if (mesh_4_6_io_out_valid_0) begin
      _T_139_0 <= mesh_4_6_io_out_b_0;
    end
    if (mesh_5_6_io_out_valid_0) begin
      _T_140_0 <= mesh_5_6_io_out_b_0;
    end
    if (mesh_6_6_io_out_valid_0) begin
      _T_141_0 <= mesh_6_6_io_out_b_0;
    end
    _T_142_0 <= io_in_d_7_0;
    _T_143_0 <= io_in_valid_7_0;
    if (_T_143_0) begin
      _T_144_0 <= _T_142_0;
    end
    if (mesh_0_7_io_out_valid_0) begin
      _T_145_0 <= mesh_0_7_io_out_b_0;
    end
    if (mesh_1_7_io_out_valid_0) begin
      _T_146_0 <= mesh_1_7_io_out_b_0;
    end
    if (mesh_2_7_io_out_valid_0) begin
      _T_147_0 <= mesh_2_7_io_out_b_0;
    end
    if (mesh_3_7_io_out_valid_0) begin
      _T_148_0 <= mesh_3_7_io_out_b_0;
    end
    if (mesh_4_7_io_out_valid_0) begin
      _T_149_0 <= mesh_4_7_io_out_b_0;
    end
    if (mesh_5_7_io_out_valid_0) begin
      _T_150_0 <= mesh_5_7_io_out_b_0;
    end
    if (mesh_6_7_io_out_valid_0) begin
      _T_151_0 <= mesh_6_7_io_out_b_0;
    end
    _T_152_0 <= io_in_b_0_0;
    _T_153_0 <= io_in_valid_0_0;
    if (_T_153_0) begin
      _T_154_0 <= _T_152_0;
    end
    if (mesh_0_0_io_out_valid_0) begin
      _T_155_0 <= mesh_0_0_io_out_c_0;
    end
    if (mesh_1_0_io_out_valid_0) begin
      _T_156_0 <= mesh_1_0_io_out_c_0;
    end
    if (mesh_2_0_io_out_valid_0) begin
      _T_157_0 <= mesh_2_0_io_out_c_0;
    end
    if (mesh_3_0_io_out_valid_0) begin
      _T_158_0 <= mesh_3_0_io_out_c_0;
    end
    if (mesh_4_0_io_out_valid_0) begin
      _T_159_0 <= mesh_4_0_io_out_c_0;
    end
    if (mesh_5_0_io_out_valid_0) begin
      _T_160_0 <= mesh_5_0_io_out_c_0;
    end
    if (mesh_6_0_io_out_valid_0) begin
      _T_161_0 <= mesh_6_0_io_out_c_0;
    end
    _T_162_0 <= io_in_b_1_0;
    _T_163_0 <= io_in_valid_1_0;
    if (_T_163_0) begin
      _T_164_0 <= _T_162_0;
    end
    if (mesh_0_1_io_out_valid_0) begin
      _T_165_0 <= mesh_0_1_io_out_c_0;
    end
    if (mesh_1_1_io_out_valid_0) begin
      _T_166_0 <= mesh_1_1_io_out_c_0;
    end
    if (mesh_2_1_io_out_valid_0) begin
      _T_167_0 <= mesh_2_1_io_out_c_0;
    end
    if (mesh_3_1_io_out_valid_0) begin
      _T_168_0 <= mesh_3_1_io_out_c_0;
    end
    if (mesh_4_1_io_out_valid_0) begin
      _T_169_0 <= mesh_4_1_io_out_c_0;
    end
    if (mesh_5_1_io_out_valid_0) begin
      _T_170_0 <= mesh_5_1_io_out_c_0;
    end
    if (mesh_6_1_io_out_valid_0) begin
      _T_171_0 <= mesh_6_1_io_out_c_0;
    end
    _T_172_0 <= io_in_b_2_0;
    _T_173_0 <= io_in_valid_2_0;
    if (_T_173_0) begin
      _T_174_0 <= _T_172_0;
    end
    if (mesh_0_2_io_out_valid_0) begin
      _T_175_0 <= mesh_0_2_io_out_c_0;
    end
    if (mesh_1_2_io_out_valid_0) begin
      _T_176_0 <= mesh_1_2_io_out_c_0;
    end
    if (mesh_2_2_io_out_valid_0) begin
      _T_177_0 <= mesh_2_2_io_out_c_0;
    end
    if (mesh_3_2_io_out_valid_0) begin
      _T_178_0 <= mesh_3_2_io_out_c_0;
    end
    if (mesh_4_2_io_out_valid_0) begin
      _T_179_0 <= mesh_4_2_io_out_c_0;
    end
    if (mesh_5_2_io_out_valid_0) begin
      _T_180_0 <= mesh_5_2_io_out_c_0;
    end
    if (mesh_6_2_io_out_valid_0) begin
      _T_181_0 <= mesh_6_2_io_out_c_0;
    end
    _T_182_0 <= io_in_b_3_0;
    _T_183_0 <= io_in_valid_3_0;
    if (_T_183_0) begin
      _T_184_0 <= _T_182_0;
    end
    if (mesh_0_3_io_out_valid_0) begin
      _T_185_0 <= mesh_0_3_io_out_c_0;
    end
    if (mesh_1_3_io_out_valid_0) begin
      _T_186_0 <= mesh_1_3_io_out_c_0;
    end
    if (mesh_2_3_io_out_valid_0) begin
      _T_187_0 <= mesh_2_3_io_out_c_0;
    end
    if (mesh_3_3_io_out_valid_0) begin
      _T_188_0 <= mesh_3_3_io_out_c_0;
    end
    if (mesh_4_3_io_out_valid_0) begin
      _T_189_0 <= mesh_4_3_io_out_c_0;
    end
    if (mesh_5_3_io_out_valid_0) begin
      _T_190_0 <= mesh_5_3_io_out_c_0;
    end
    if (mesh_6_3_io_out_valid_0) begin
      _T_191_0 <= mesh_6_3_io_out_c_0;
    end
    _T_192_0 <= io_in_b_4_0;
    _T_193_0 <= io_in_valid_4_0;
    if (_T_193_0) begin
      _T_194_0 <= _T_192_0;
    end
    if (mesh_0_4_io_out_valid_0) begin
      _T_195_0 <= mesh_0_4_io_out_c_0;
    end
    if (mesh_1_4_io_out_valid_0) begin
      _T_196_0 <= mesh_1_4_io_out_c_0;
    end
    if (mesh_2_4_io_out_valid_0) begin
      _T_197_0 <= mesh_2_4_io_out_c_0;
    end
    if (mesh_3_4_io_out_valid_0) begin
      _T_198_0 <= mesh_3_4_io_out_c_0;
    end
    if (mesh_4_4_io_out_valid_0) begin
      _T_199_0 <= mesh_4_4_io_out_c_0;
    end
    if (mesh_5_4_io_out_valid_0) begin
      _T_200_0 <= mesh_5_4_io_out_c_0;
    end
    if (mesh_6_4_io_out_valid_0) begin
      _T_201_0 <= mesh_6_4_io_out_c_0;
    end
    _T_202_0 <= io_in_b_5_0;
    _T_203_0 <= io_in_valid_5_0;
    if (_T_203_0) begin
      _T_204_0 <= _T_202_0;
    end
    if (mesh_0_5_io_out_valid_0) begin
      _T_205_0 <= mesh_0_5_io_out_c_0;
    end
    if (mesh_1_5_io_out_valid_0) begin
      _T_206_0 <= mesh_1_5_io_out_c_0;
    end
    if (mesh_2_5_io_out_valid_0) begin
      _T_207_0 <= mesh_2_5_io_out_c_0;
    end
    if (mesh_3_5_io_out_valid_0) begin
      _T_208_0 <= mesh_3_5_io_out_c_0;
    end
    if (mesh_4_5_io_out_valid_0) begin
      _T_209_0 <= mesh_4_5_io_out_c_0;
    end
    if (mesh_5_5_io_out_valid_0) begin
      _T_210_0 <= mesh_5_5_io_out_c_0;
    end
    if (mesh_6_5_io_out_valid_0) begin
      _T_211_0 <= mesh_6_5_io_out_c_0;
    end
    _T_212_0 <= io_in_b_6_0;
    _T_213_0 <= io_in_valid_6_0;
    if (_T_213_0) begin
      _T_214_0 <= _T_212_0;
    end
    if (mesh_0_6_io_out_valid_0) begin
      _T_215_0 <= mesh_0_6_io_out_c_0;
    end
    if (mesh_1_6_io_out_valid_0) begin
      _T_216_0 <= mesh_1_6_io_out_c_0;
    end
    if (mesh_2_6_io_out_valid_0) begin
      _T_217_0 <= mesh_2_6_io_out_c_0;
    end
    if (mesh_3_6_io_out_valid_0) begin
      _T_218_0 <= mesh_3_6_io_out_c_0;
    end
    if (mesh_4_6_io_out_valid_0) begin
      _T_219_0 <= mesh_4_6_io_out_c_0;
    end
    if (mesh_5_6_io_out_valid_0) begin
      _T_220_0 <= mesh_5_6_io_out_c_0;
    end
    if (mesh_6_6_io_out_valid_0) begin
      _T_221_0 <= mesh_6_6_io_out_c_0;
    end
    _T_222_0 <= io_in_b_7_0;
    _T_223_0 <= io_in_valid_7_0;
    if (_T_223_0) begin
      _T_224_0 <= _T_222_0;
    end
    if (mesh_0_7_io_out_valid_0) begin
      _T_225_0 <= mesh_0_7_io_out_c_0;
    end
    if (mesh_1_7_io_out_valid_0) begin
      _T_226_0 <= mesh_1_7_io_out_c_0;
    end
    if (mesh_2_7_io_out_valid_0) begin
      _T_227_0 <= mesh_2_7_io_out_c_0;
    end
    if (mesh_3_7_io_out_valid_0) begin
      _T_228_0 <= mesh_3_7_io_out_c_0;
    end
    if (mesh_4_7_io_out_valid_0) begin
      _T_229_0 <= mesh_4_7_io_out_c_0;
    end
    if (mesh_5_7_io_out_valid_0) begin
      _T_230_0 <= mesh_5_7_io_out_c_0;
    end
    if (mesh_6_7_io_out_valid_0) begin
      _T_231_0 <= mesh_6_7_io_out_c_0;
    end
    _T_232_0_propagate <= io_in_control_0_0_propagate;
    _T_232_0_shift <= io_in_control_0_0_shift;
    _T_233_0 <= io_in_valid_0_0;
    if (_T_233_0) begin
      _T_234 <= _T_232_0_shift;
    end
    if (_T_233_0) begin
      _T_236 <= _T_232_0_propagate;
    end
    if (mesh_0_0_io_out_valid_0) begin
      _T_237 <= mesh_0_0_io_out_control_0_shift;
    end
    if (mesh_0_0_io_out_valid_0) begin
      _T_239 <= mesh_0_0_io_out_control_0_propagate;
    end
    if (mesh_1_0_io_out_valid_0) begin
      _T_240 <= mesh_1_0_io_out_control_0_shift;
    end
    if (mesh_1_0_io_out_valid_0) begin
      _T_242 <= mesh_1_0_io_out_control_0_propagate;
    end
    if (mesh_2_0_io_out_valid_0) begin
      _T_243 <= mesh_2_0_io_out_control_0_shift;
    end
    if (mesh_2_0_io_out_valid_0) begin
      _T_245 <= mesh_2_0_io_out_control_0_propagate;
    end
    if (mesh_3_0_io_out_valid_0) begin
      _T_246 <= mesh_3_0_io_out_control_0_shift;
    end
    if (mesh_3_0_io_out_valid_0) begin
      _T_248 <= mesh_3_0_io_out_control_0_propagate;
    end
    if (mesh_4_0_io_out_valid_0) begin
      _T_249 <= mesh_4_0_io_out_control_0_shift;
    end
    if (mesh_4_0_io_out_valid_0) begin
      _T_251 <= mesh_4_0_io_out_control_0_propagate;
    end
    if (mesh_5_0_io_out_valid_0) begin
      _T_252 <= mesh_5_0_io_out_control_0_shift;
    end
    if (mesh_5_0_io_out_valid_0) begin
      _T_254 <= mesh_5_0_io_out_control_0_propagate;
    end
    if (mesh_6_0_io_out_valid_0) begin
      _T_255 <= mesh_6_0_io_out_control_0_shift;
    end
    if (mesh_6_0_io_out_valid_0) begin
      _T_257 <= mesh_6_0_io_out_control_0_propagate;
    end
    _T_258_0_propagate <= io_in_control_1_0_propagate;
    _T_258_0_shift <= io_in_control_1_0_shift;
    _T_259_0 <= io_in_valid_1_0;
    if (_T_259_0) begin
      _T_260 <= _T_258_0_shift;
    end
    if (_T_259_0) begin
      _T_262 <= _T_258_0_propagate;
    end
    if (mesh_0_1_io_out_valid_0) begin
      _T_263 <= mesh_0_1_io_out_control_0_shift;
    end
    if (mesh_0_1_io_out_valid_0) begin
      _T_265 <= mesh_0_1_io_out_control_0_propagate;
    end
    if (mesh_1_1_io_out_valid_0) begin
      _T_266 <= mesh_1_1_io_out_control_0_shift;
    end
    if (mesh_1_1_io_out_valid_0) begin
      _T_268 <= mesh_1_1_io_out_control_0_propagate;
    end
    if (mesh_2_1_io_out_valid_0) begin
      _T_269 <= mesh_2_1_io_out_control_0_shift;
    end
    if (mesh_2_1_io_out_valid_0) begin
      _T_271 <= mesh_2_1_io_out_control_0_propagate;
    end
    if (mesh_3_1_io_out_valid_0) begin
      _T_272 <= mesh_3_1_io_out_control_0_shift;
    end
    if (mesh_3_1_io_out_valid_0) begin
      _T_274 <= mesh_3_1_io_out_control_0_propagate;
    end
    if (mesh_4_1_io_out_valid_0) begin
      _T_275 <= mesh_4_1_io_out_control_0_shift;
    end
    if (mesh_4_1_io_out_valid_0) begin
      _T_277 <= mesh_4_1_io_out_control_0_propagate;
    end
    if (mesh_5_1_io_out_valid_0) begin
      _T_278 <= mesh_5_1_io_out_control_0_shift;
    end
    if (mesh_5_1_io_out_valid_0) begin
      _T_280 <= mesh_5_1_io_out_control_0_propagate;
    end
    if (mesh_6_1_io_out_valid_0) begin
      _T_281 <= mesh_6_1_io_out_control_0_shift;
    end
    if (mesh_6_1_io_out_valid_0) begin
      _T_283 <= mesh_6_1_io_out_control_0_propagate;
    end
    _T_284_0_propagate <= io_in_control_2_0_propagate;
    _T_284_0_shift <= io_in_control_2_0_shift;
    _T_285_0 <= io_in_valid_2_0;
    if (_T_285_0) begin
      _T_286 <= _T_284_0_shift;
    end
    if (_T_285_0) begin
      _T_288 <= _T_284_0_propagate;
    end
    if (mesh_0_2_io_out_valid_0) begin
      _T_289 <= mesh_0_2_io_out_control_0_shift;
    end
    if (mesh_0_2_io_out_valid_0) begin
      _T_291 <= mesh_0_2_io_out_control_0_propagate;
    end
    if (mesh_1_2_io_out_valid_0) begin
      _T_292 <= mesh_1_2_io_out_control_0_shift;
    end
    if (mesh_1_2_io_out_valid_0) begin
      _T_294 <= mesh_1_2_io_out_control_0_propagate;
    end
    if (mesh_2_2_io_out_valid_0) begin
      _T_295 <= mesh_2_2_io_out_control_0_shift;
    end
    if (mesh_2_2_io_out_valid_0) begin
      _T_297 <= mesh_2_2_io_out_control_0_propagate;
    end
    if (mesh_3_2_io_out_valid_0) begin
      _T_298 <= mesh_3_2_io_out_control_0_shift;
    end
    if (mesh_3_2_io_out_valid_0) begin
      _T_300 <= mesh_3_2_io_out_control_0_propagate;
    end
    if (mesh_4_2_io_out_valid_0) begin
      _T_301 <= mesh_4_2_io_out_control_0_shift;
    end
    if (mesh_4_2_io_out_valid_0) begin
      _T_303 <= mesh_4_2_io_out_control_0_propagate;
    end
    if (mesh_5_2_io_out_valid_0) begin
      _T_304 <= mesh_5_2_io_out_control_0_shift;
    end
    if (mesh_5_2_io_out_valid_0) begin
      _T_306 <= mesh_5_2_io_out_control_0_propagate;
    end
    if (mesh_6_2_io_out_valid_0) begin
      _T_307 <= mesh_6_2_io_out_control_0_shift;
    end
    if (mesh_6_2_io_out_valid_0) begin
      _T_309 <= mesh_6_2_io_out_control_0_propagate;
    end
    _T_310_0_propagate <= io_in_control_3_0_propagate;
    _T_310_0_shift <= io_in_control_3_0_shift;
    _T_311_0 <= io_in_valid_3_0;
    if (_T_311_0) begin
      _T_312 <= _T_310_0_shift;
    end
    if (_T_311_0) begin
      _T_314 <= _T_310_0_propagate;
    end
    if (mesh_0_3_io_out_valid_0) begin
      _T_315 <= mesh_0_3_io_out_control_0_shift;
    end
    if (mesh_0_3_io_out_valid_0) begin
      _T_317 <= mesh_0_3_io_out_control_0_propagate;
    end
    if (mesh_1_3_io_out_valid_0) begin
      _T_318 <= mesh_1_3_io_out_control_0_shift;
    end
    if (mesh_1_3_io_out_valid_0) begin
      _T_320 <= mesh_1_3_io_out_control_0_propagate;
    end
    if (mesh_2_3_io_out_valid_0) begin
      _T_321 <= mesh_2_3_io_out_control_0_shift;
    end
    if (mesh_2_3_io_out_valid_0) begin
      _T_323 <= mesh_2_3_io_out_control_0_propagate;
    end
    if (mesh_3_3_io_out_valid_0) begin
      _T_324 <= mesh_3_3_io_out_control_0_shift;
    end
    if (mesh_3_3_io_out_valid_0) begin
      _T_326 <= mesh_3_3_io_out_control_0_propagate;
    end
    if (mesh_4_3_io_out_valid_0) begin
      _T_327 <= mesh_4_3_io_out_control_0_shift;
    end
    if (mesh_4_3_io_out_valid_0) begin
      _T_329 <= mesh_4_3_io_out_control_0_propagate;
    end
    if (mesh_5_3_io_out_valid_0) begin
      _T_330 <= mesh_5_3_io_out_control_0_shift;
    end
    if (mesh_5_3_io_out_valid_0) begin
      _T_332 <= mesh_5_3_io_out_control_0_propagate;
    end
    if (mesh_6_3_io_out_valid_0) begin
      _T_333 <= mesh_6_3_io_out_control_0_shift;
    end
    if (mesh_6_3_io_out_valid_0) begin
      _T_335 <= mesh_6_3_io_out_control_0_propagate;
    end
    _T_336_0_propagate <= io_in_control_4_0_propagate;
    _T_336_0_shift <= io_in_control_4_0_shift;
    _T_337_0 <= io_in_valid_4_0;
    if (_T_337_0) begin
      _T_338 <= _T_336_0_shift;
    end
    if (_T_337_0) begin
      _T_340 <= _T_336_0_propagate;
    end
    if (mesh_0_4_io_out_valid_0) begin
      _T_341 <= mesh_0_4_io_out_control_0_shift;
    end
    if (mesh_0_4_io_out_valid_0) begin
      _T_343 <= mesh_0_4_io_out_control_0_propagate;
    end
    if (mesh_1_4_io_out_valid_0) begin
      _T_344 <= mesh_1_4_io_out_control_0_shift;
    end
    if (mesh_1_4_io_out_valid_0) begin
      _T_346 <= mesh_1_4_io_out_control_0_propagate;
    end
    if (mesh_2_4_io_out_valid_0) begin
      _T_347 <= mesh_2_4_io_out_control_0_shift;
    end
    if (mesh_2_4_io_out_valid_0) begin
      _T_349 <= mesh_2_4_io_out_control_0_propagate;
    end
    if (mesh_3_4_io_out_valid_0) begin
      _T_350 <= mesh_3_4_io_out_control_0_shift;
    end
    if (mesh_3_4_io_out_valid_0) begin
      _T_352 <= mesh_3_4_io_out_control_0_propagate;
    end
    if (mesh_4_4_io_out_valid_0) begin
      _T_353 <= mesh_4_4_io_out_control_0_shift;
    end
    if (mesh_4_4_io_out_valid_0) begin
      _T_355 <= mesh_4_4_io_out_control_0_propagate;
    end
    if (mesh_5_4_io_out_valid_0) begin
      _T_356 <= mesh_5_4_io_out_control_0_shift;
    end
    if (mesh_5_4_io_out_valid_0) begin
      _T_358 <= mesh_5_4_io_out_control_0_propagate;
    end
    if (mesh_6_4_io_out_valid_0) begin
      _T_359 <= mesh_6_4_io_out_control_0_shift;
    end
    if (mesh_6_4_io_out_valid_0) begin
      _T_361 <= mesh_6_4_io_out_control_0_propagate;
    end
    _T_362_0_propagate <= io_in_control_5_0_propagate;
    _T_362_0_shift <= io_in_control_5_0_shift;
    _T_363_0 <= io_in_valid_5_0;
    if (_T_363_0) begin
      _T_364 <= _T_362_0_shift;
    end
    if (_T_363_0) begin
      _T_366 <= _T_362_0_propagate;
    end
    if (mesh_0_5_io_out_valid_0) begin
      _T_367 <= mesh_0_5_io_out_control_0_shift;
    end
    if (mesh_0_5_io_out_valid_0) begin
      _T_369 <= mesh_0_5_io_out_control_0_propagate;
    end
    if (mesh_1_5_io_out_valid_0) begin
      _T_370 <= mesh_1_5_io_out_control_0_shift;
    end
    if (mesh_1_5_io_out_valid_0) begin
      _T_372 <= mesh_1_5_io_out_control_0_propagate;
    end
    if (mesh_2_5_io_out_valid_0) begin
      _T_373 <= mesh_2_5_io_out_control_0_shift;
    end
    if (mesh_2_5_io_out_valid_0) begin
      _T_375 <= mesh_2_5_io_out_control_0_propagate;
    end
    if (mesh_3_5_io_out_valid_0) begin
      _T_376 <= mesh_3_5_io_out_control_0_shift;
    end
    if (mesh_3_5_io_out_valid_0) begin
      _T_378 <= mesh_3_5_io_out_control_0_propagate;
    end
    if (mesh_4_5_io_out_valid_0) begin
      _T_379 <= mesh_4_5_io_out_control_0_shift;
    end
    if (mesh_4_5_io_out_valid_0) begin
      _T_381 <= mesh_4_5_io_out_control_0_propagate;
    end
    if (mesh_5_5_io_out_valid_0) begin
      _T_382 <= mesh_5_5_io_out_control_0_shift;
    end
    if (mesh_5_5_io_out_valid_0) begin
      _T_384 <= mesh_5_5_io_out_control_0_propagate;
    end
    if (mesh_6_5_io_out_valid_0) begin
      _T_385 <= mesh_6_5_io_out_control_0_shift;
    end
    if (mesh_6_5_io_out_valid_0) begin
      _T_387 <= mesh_6_5_io_out_control_0_propagate;
    end
    _T_388_0_propagate <= io_in_control_6_0_propagate;
    _T_388_0_shift <= io_in_control_6_0_shift;
    _T_389_0 <= io_in_valid_6_0;
    if (_T_389_0) begin
      _T_390 <= _T_388_0_shift;
    end
    if (_T_389_0) begin
      _T_392 <= _T_388_0_propagate;
    end
    if (mesh_0_6_io_out_valid_0) begin
      _T_393 <= mesh_0_6_io_out_control_0_shift;
    end
    if (mesh_0_6_io_out_valid_0) begin
      _T_395 <= mesh_0_6_io_out_control_0_propagate;
    end
    if (mesh_1_6_io_out_valid_0) begin
      _T_396 <= mesh_1_6_io_out_control_0_shift;
    end
    if (mesh_1_6_io_out_valid_0) begin
      _T_398 <= mesh_1_6_io_out_control_0_propagate;
    end
    if (mesh_2_6_io_out_valid_0) begin
      _T_399 <= mesh_2_6_io_out_control_0_shift;
    end
    if (mesh_2_6_io_out_valid_0) begin
      _T_401 <= mesh_2_6_io_out_control_0_propagate;
    end
    if (mesh_3_6_io_out_valid_0) begin
      _T_402 <= mesh_3_6_io_out_control_0_shift;
    end
    if (mesh_3_6_io_out_valid_0) begin
      _T_404 <= mesh_3_6_io_out_control_0_propagate;
    end
    if (mesh_4_6_io_out_valid_0) begin
      _T_405 <= mesh_4_6_io_out_control_0_shift;
    end
    if (mesh_4_6_io_out_valid_0) begin
      _T_407 <= mesh_4_6_io_out_control_0_propagate;
    end
    if (mesh_5_6_io_out_valid_0) begin
      _T_408 <= mesh_5_6_io_out_control_0_shift;
    end
    if (mesh_5_6_io_out_valid_0) begin
      _T_410 <= mesh_5_6_io_out_control_0_propagate;
    end
    if (mesh_6_6_io_out_valid_0) begin
      _T_411 <= mesh_6_6_io_out_control_0_shift;
    end
    if (mesh_6_6_io_out_valid_0) begin
      _T_413 <= mesh_6_6_io_out_control_0_propagate;
    end
    _T_414_0_propagate <= io_in_control_7_0_propagate;
    _T_414_0_shift <= io_in_control_7_0_shift;
    _T_415_0 <= io_in_valid_7_0;
    if (_T_415_0) begin
      _T_416 <= _T_414_0_shift;
    end
    if (_T_415_0) begin
      _T_418 <= _T_414_0_propagate;
    end
    if (mesh_0_7_io_out_valid_0) begin
      _T_419 <= mesh_0_7_io_out_control_0_shift;
    end
    if (mesh_0_7_io_out_valid_0) begin
      _T_421 <= mesh_0_7_io_out_control_0_propagate;
    end
    if (mesh_1_7_io_out_valid_0) begin
      _T_422 <= mesh_1_7_io_out_control_0_shift;
    end
    if (mesh_1_7_io_out_valid_0) begin
      _T_424 <= mesh_1_7_io_out_control_0_propagate;
    end
    if (mesh_2_7_io_out_valid_0) begin
      _T_425 <= mesh_2_7_io_out_control_0_shift;
    end
    if (mesh_2_7_io_out_valid_0) begin
      _T_427 <= mesh_2_7_io_out_control_0_propagate;
    end
    if (mesh_3_7_io_out_valid_0) begin
      _T_428 <= mesh_3_7_io_out_control_0_shift;
    end
    if (mesh_3_7_io_out_valid_0) begin
      _T_430 <= mesh_3_7_io_out_control_0_propagate;
    end
    if (mesh_4_7_io_out_valid_0) begin
      _T_431 <= mesh_4_7_io_out_control_0_shift;
    end
    if (mesh_4_7_io_out_valid_0) begin
      _T_433 <= mesh_4_7_io_out_control_0_propagate;
    end
    if (mesh_5_7_io_out_valid_0) begin
      _T_434 <= mesh_5_7_io_out_control_0_shift;
    end
    if (mesh_5_7_io_out_valid_0) begin
      _T_436 <= mesh_5_7_io_out_control_0_propagate;
    end
    if (mesh_6_7_io_out_valid_0) begin
      _T_437 <= mesh_6_7_io_out_control_0_shift;
    end
    if (mesh_6_7_io_out_valid_0) begin
      _T_439 <= mesh_6_7_io_out_control_0_propagate;
    end
    _T_440_0 <= io_in_valid_0_0;
    _T_441_0 <= _T_440_0;
    _T_442_0 <= mesh_0_0_io_out_valid_0;
    _T_443_0 <= mesh_1_0_io_out_valid_0;
    _T_444_0 <= mesh_2_0_io_out_valid_0;
    _T_445_0 <= mesh_3_0_io_out_valid_0;
    _T_446_0 <= mesh_4_0_io_out_valid_0;
    _T_447_0 <= mesh_5_0_io_out_valid_0;
    _T_448_0 <= mesh_6_0_io_out_valid_0;
    _T_449_0 <= io_in_valid_1_0;
    _T_450_0 <= _T_449_0;
    _T_451_0 <= mesh_0_1_io_out_valid_0;
    _T_452_0 <= mesh_1_1_io_out_valid_0;
    _T_453_0 <= mesh_2_1_io_out_valid_0;
    _T_454_0 <= mesh_3_1_io_out_valid_0;
    _T_455_0 <= mesh_4_1_io_out_valid_0;
    _T_456_0 <= mesh_5_1_io_out_valid_0;
    _T_457_0 <= mesh_6_1_io_out_valid_0;
    _T_458_0 <= io_in_valid_2_0;
    _T_459_0 <= _T_458_0;
    _T_460_0 <= mesh_0_2_io_out_valid_0;
    _T_461_0 <= mesh_1_2_io_out_valid_0;
    _T_462_0 <= mesh_2_2_io_out_valid_0;
    _T_463_0 <= mesh_3_2_io_out_valid_0;
    _T_464_0 <= mesh_4_2_io_out_valid_0;
    _T_465_0 <= mesh_5_2_io_out_valid_0;
    _T_466_0 <= mesh_6_2_io_out_valid_0;
    _T_467_0 <= io_in_valid_3_0;
    _T_468_0 <= _T_467_0;
    _T_469_0 <= mesh_0_3_io_out_valid_0;
    _T_470_0 <= mesh_1_3_io_out_valid_0;
    _T_471_0 <= mesh_2_3_io_out_valid_0;
    _T_472_0 <= mesh_3_3_io_out_valid_0;
    _T_473_0 <= mesh_4_3_io_out_valid_0;
    _T_474_0 <= mesh_5_3_io_out_valid_0;
    _T_475_0 <= mesh_6_3_io_out_valid_0;
    _T_476_0 <= io_in_valid_4_0;
    _T_477_0 <= _T_476_0;
    _T_478_0 <= mesh_0_4_io_out_valid_0;
    _T_479_0 <= mesh_1_4_io_out_valid_0;
    _T_480_0 <= mesh_2_4_io_out_valid_0;
    _T_481_0 <= mesh_3_4_io_out_valid_0;
    _T_482_0 <= mesh_4_4_io_out_valid_0;
    _T_483_0 <= mesh_5_4_io_out_valid_0;
    _T_484_0 <= mesh_6_4_io_out_valid_0;
    _T_485_0 <= io_in_valid_5_0;
    _T_486_0 <= _T_485_0;
    _T_487_0 <= mesh_0_5_io_out_valid_0;
    _T_488_0 <= mesh_1_5_io_out_valid_0;
    _T_489_0 <= mesh_2_5_io_out_valid_0;
    _T_490_0 <= mesh_3_5_io_out_valid_0;
    _T_491_0 <= mesh_4_5_io_out_valid_0;
    _T_492_0 <= mesh_5_5_io_out_valid_0;
    _T_493_0 <= mesh_6_5_io_out_valid_0;
    _T_494_0 <= io_in_valid_6_0;
    _T_495_0 <= _T_494_0;
    _T_496_0 <= mesh_0_6_io_out_valid_0;
    _T_497_0 <= mesh_1_6_io_out_valid_0;
    _T_498_0 <= mesh_2_6_io_out_valid_0;
    _T_499_0 <= mesh_3_6_io_out_valid_0;
    _T_500_0 <= mesh_4_6_io_out_valid_0;
    _T_501_0 <= mesh_5_6_io_out_valid_0;
    _T_502_0 <= mesh_6_6_io_out_valid_0;
    _T_503_0 <= io_in_valid_7_0;
    _T_504_0 <= _T_503_0;
    _T_505_0 <= mesh_0_7_io_out_valid_0;
    _T_506_0 <= mesh_1_7_io_out_valid_0;
    _T_507_0 <= mesh_2_7_io_out_valid_0;
    _T_508_0 <= mesh_3_7_io_out_valid_0;
    _T_509_0 <= mesh_4_7_io_out_valid_0;
    _T_510_0 <= mesh_5_7_io_out_valid_0;
    _T_511_0 <= mesh_6_7_io_out_valid_0;
  end
endmodule
